
//
// Verific Verilog Description of module top
//

module top (clk, clk_0, clk_1, o_pllBr0_reg, o_pllBr1_reg, bscan_DRCK, 
            bscan_RESET, bscan_TMS, bscan_RUNTEST, bscan_SEL, bscan_SHIFT, 
            bscan_TDI, bscan_CAPTURE, bscan_TCK, bscan_UPDATE, bscan_TDO);
    input clk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/top.v(2)
    input clk_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/top.v(4)
    input clk_1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/top.v(5)
    output [255:0]o_pllBr0_reg /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/top.v(7)
    output [255:0]o_pllBr1_reg /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/top.v(8)
    input bscan_DRCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/top.v(10)
    input bscan_RESET /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/top.v(11)
    input bscan_TMS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/top.v(12)
    input bscan_RUNTEST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/top.v(13)
    input bscan_SEL /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/top.v(14)
    input bscan_SHIFT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/top.v(15)
    input bscan_TDI /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/top.v(16)
    input bscan_CAPTURE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/top.v(17)
    input bscan_TCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/top.v(18)
    input bscan_UPDATE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/top.v(19)
    output bscan_TDO /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/top.v(20)
    
    wire [255:0]\test_module/n33 ;
    
    wire \test_module/add_41/n180 , \test_module/add_41/n172 , \test_module/add_41/n190 , 
        \test_module/add_41/n2 , \test_module/add_41/n170 ;
    wire [20:0]\test_module/n1132 ;
    
    wire \test_module/add_44/n2 , \test_module/add_41/n192 ;
    wire [20:0]\test_module/delay_1 ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(10)
    
    wire \test_module/add_41/n168 , \test_module/add_41/n166 ;
    wire [255:0]\test_module/n1156 ;
    
    wire \test_module/add_46/n2 ;
    wire [5:0]\debug_inst/vio0/vio_core_inst/n408 ;
    
    wire \debug_inst/vio0/vio_core_inst/add_772/n2 , \test_module/add_41/n194 ;
    wire [20:0]\test_module/delay_2 ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(10)
    
    wire \test_module/add_41/n164 , \test_module/add_41/n162 , \test_module/add_41/n160 , 
        \test_module/add_41/n158 , \test_module/add_41/n156 , \test_module/add_41/n154 , 
        \test_module/add_41/n152 , \test_module/add_41/n150 , \test_module/add_41/n148 , 
        \test_module/add_41/n196 , \test_module/add_41/n198 , \test_module/add_41/n200 , 
        \test_module/add_41/n202 , \test_module/add_41/n204 , \test_module/add_41/n206 , 
        \test_module/add_41/n208 , \test_module/add_41/n210 , \test_module/add_41/n212 , 
        \test_module/add_41/n214 , \test_module/add_41/n216 , \test_module/add_41/n218 , 
        \test_module/add_41/n220 , \test_module/add_41/n222 , \test_module/add_41/n224 , 
        \test_module/add_41/n226 , \test_module/add_41/n228 , \test_module/add_41/n230 , 
        \test_module/add_41/n232 , \test_module/add_41/n234 , \test_module/add_41/n236 , 
        \test_module/add_41/n146 , \test_module/add_41/n144 , \test_module/add_41/n142 , 
        \test_module/add_41/n140 , \test_module/add_41/n138 , \test_module/add_41/n136 , 
        \test_module/add_41/n134 , \test_module/add_41/n238 , \test_module/add_41/n240 , 
        \test_module/add_41/n242 , \test_module/add_41/n244 , \test_module/add_41/n246 , 
        \test_module/add_41/n248 , \test_module/add_41/n250 , \test_module/add_41/n252 , 
        \test_module/add_41/n254 , \test_module/add_41/n256 , \test_module/add_41/n258 , 
        \test_module/add_41/n260 , \test_module/add_41/n262 , \test_module/add_41/n264 , 
        \test_module/add_41/n266 , \test_module/add_41/n268 , \test_module/add_41/n270 , 
        \test_module/add_41/n272 , \test_module/add_41/n274 , \test_module/add_41/n276 , 
        \test_module/add_41/n278 ;
    wire [2:0]\debug_inst/vio0/vio_core_inst/internal_reg_r0 ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1185)
    wire [32:0]\debug_inst/vio0/vio_core_inst/incremented_address ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1237)
    
    wire \debug_inst/vio0/vio_core_inst/add_33/n4 ;
    wire [5:0]\debug_inst/vio0/vio_core_inst/bit_count ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1190)
    
    wire \test_module/add_41/n132 , \test_module/add_41/n130 , \test_module/add_41/n178 , 
        \test_module/add_41/n184 , \test_module/add_41/n280 , \test_module/add_41/n282 ;
    wire [15:0]\debug_inst/vio0/vio_core_inst/word_count ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1191)
    wire [15:0]\debug_inst/vio0/vio_core_inst/data_out_shift_reg ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1186)
    
    wire \test_module/add_41/n284 ;
    wire [3:0]\debug_inst/vio0/vio_core_inst/module_state ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1246)
    
    wire \test_module/add_41/n176 ;
    wire [15:0]\debug_inst/vio0/vio_core_inst/data_from_biu ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1244)
    
    wire \test_module/add_41/n128 , \test_module/add_41/n126 , \test_module/add_41/n124 , 
        \test_module/add_41/n122 , \test_module/add_41/n120 , \test_module/add_41/n118 , 
        \test_module/add_41/n116 , \test_module/add_41/n114 , \test_module/add_41/n112 , 
        \test_module/add_41/n110 , \test_module/add_41/n108 , \test_module/add_41/n106 , 
        \test_module/add_41/n104 , \test_module/add_41/n102 , \test_module/add_41/n286 , 
        \test_module/add_41/n288 , \test_module/add_41/n290 , \test_module/add_41/n292 , 
        \test_module/add_41/n294 , \test_module/add_41/n296 , \test_module/add_41/n298 , 
        \test_module/add_41/n300 , \test_module/add_41/n302 , \test_module/add_41/n304 , 
        \test_module/add_41/n306 , \test_module/add_41/n308 , \test_module/add_41/n310 , 
        \test_module/add_41/n312 , \test_module/add_41/n314 , \test_module/add_41/n316 , 
        \test_module/add_41/n318 , \test_module/add_41/n320 , \test_module/add_41/n322 , 
        \test_module/add_41/n324 , \test_module/add_41/n326 , \test_module/add_41/n328 , 
        \test_module/add_41/n330 , \test_module/add_41/n332 , \test_module/add_41/n334 , 
        \test_module/add_41/n336 , \test_module/add_41/n338 , \test_module/add_41/n340 , 
        \test_module/add_41/n342 , \test_module/add_41/n344 , \test_module/add_41/n346 , 
        \test_module/add_41/n348 , \test_module/add_41/n350 , \test_module/add_41/n352 , 
        \test_module/add_41/n354 , \test_module/add_41/n356 , \test_module/add_41/n358 , 
        \test_module/add_41/n360 , \test_module/add_41/n362 , \test_module/add_41/n364 , 
        \test_module/add_41/n366 , \test_module/add_41/n368 , \test_module/add_41/n370 , 
        \test_module/add_41/n372 , \test_module/add_41/n374 , \test_module/add_41/n376 , 
        \test_module/add_41/n378 , \test_module/add_41/n380 , \test_module/add_41/n382 , 
        \test_module/add_41/n384 , \test_module/add_41/n386 , \test_module/add_41/n388 , 
        \test_module/add_41/n390 , \test_module/add_41/n392 , \test_module/add_41/n394 , 
        \test_module/add_41/n396 , \test_module/add_41/n398 , \test_module/add_41/n400 , 
        \test_module/add_41/n402 , \test_module/add_41/n404 , \test_module/add_41/n406 , 
        \test_module/add_41/n408 , \test_module/add_41/n410 , \test_module/add_41/n412 , 
        \test_module/add_41/n414 , \test_module/add_41/n416 , \test_module/add_41/n418 , 
        \test_module/add_41/n420 , \test_module/add_41/n422 , \test_module/add_41/n424 , 
        \test_module/add_41/n426 ;
    wire [31:0]\debug_inst/vio0/vio_core_inst/crc_data_out ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1242)
    
    wire \test_module/add_41/n428 , \test_module/add_41/n430 , \test_module/add_41/n432 , 
        \test_module/add_41/n434 , \test_module/add_41/n436 , \test_module/add_41/n438 , 
        \test_module/add_41/n440 , \test_module/add_41/n442 , \test_module/add_41/n444 , 
        \test_module/add_41/n446 , \test_module/add_41/n448 , \test_module/add_41/n450 , 
        \test_module/add_41/n452 , \test_module/add_41/n454 , \test_module/add_41/n456 , 
        \test_module/add_41/n458 , \test_module/add_41/n460 , \test_module/add_41/n462 , 
        \test_module/add_41/n464 , \test_module/add_41/n466 , \test_module/add_41/n468 , 
        \test_module/add_41/n470 , \test_module/add_41/n472 , \test_module/add_41/n474 , 
        \test_module/add_41/n476 , \test_module/add_41/n478 , \test_module/add_41/n480 , 
        \test_module/add_41/n482 , \test_module/add_41/n484 , \test_module/add_41/n486 , 
        \test_module/add_41/n488 , \test_module/add_41/n490 , \test_module/add_41/n492 , 
        \test_module/add_41/n494 , \test_module/add_41/n496 , \test_module/add_41/n498 , 
        \test_module/add_41/n500 , \test_module/add_41/n502 , \test_module/add_41/n504 , 
        \test_module/add_41/n506 , \test_module/add_41/n508 , \test_module/add_44/n4 , 
        \test_module/add_44/n6 , \test_module/add_44/n8 , \test_module/add_44/n10 , 
        \test_module/add_44/n12 , \test_module/add_44/n14 , \test_module/add_44/n16 , 
        \test_module/add_44/n18 , \test_module/add_44/n20 , \test_module/add_44/n22 , 
        \test_module/add_44/n24 , \test_module/add_46/n4 , \test_module/add_46/n6 , 
        \test_module/add_46/n8 , \test_module/add_46/n10 , \test_module/add_46/n12 , 
        \test_module/add_46/n14 , \test_module/add_46/n16 , \test_module/add_46/n18 , 
        \test_module/add_46/n20 , \test_module/add_46/n22 , \test_module/add_46/n24 , 
        \test_module/add_46/n26 , \test_module/add_46/n28 , \test_module/add_46/n30 , 
        \test_module/add_46/n32 , \test_module/add_46/n34 , \test_module/add_46/n36 , 
        \test_module/add_46/n38 , \test_module/add_46/n40 , \test_module/add_46/n42 , 
        \test_module/add_46/n44 , \test_module/add_46/n46 , \test_module/add_46/n48 , 
        \test_module/add_46/n50 , \test_module/add_46/n52 , \test_module/add_46/n54 , 
        \test_module/add_46/n56 , \test_module/add_46/n58 , \test_module/add_46/n60 , 
        \test_module/add_46/n62 , \test_module/add_46/n64 , \test_module/add_46/n66 , 
        \test_module/add_46/n68 , \test_module/add_46/n70 , \test_module/add_46/n72 , 
        \test_module/add_46/n74 , \test_module/add_46/n76 , \test_module/add_46/n78 , 
        \test_module/add_46/n80 , \test_module/add_46/n82 , \test_module/add_46/n84 , 
        \test_module/add_46/n86 , \test_module/add_46/n88 , \test_module/add_46/n90 , 
        \test_module/add_46/n92 , \test_module/add_46/n94 , \test_module/add_46/n96 , 
        \test_module/add_46/n98 , \test_module/add_46/n100 , \test_module/add_46/n102 , 
        \test_module/add_46/n104 , \test_module/add_46/n106 , \test_module/add_46/n108 , 
        \test_module/add_46/n110 , \test_module/add_46/n112 , \test_module/add_46/n114 , 
        \test_module/add_46/n116 , \test_module/add_46/n118 , \test_module/add_46/n120 , 
        \test_module/add_46/n122 , \test_module/add_46/n124 , \test_module/add_46/n126 , 
        \test_module/add_46/n128 , \test_module/add_46/n130 , \test_module/add_46/n132 , 
        \test_module/add_46/n134 , \test_module/add_46/n136 , \test_module/add_46/n138 , 
        \test_module/add_46/n140 , \test_module/add_46/n142 , \test_module/add_46/n144 , 
        \test_module/add_46/n146 , \test_module/add_46/n148 , \test_module/add_46/n150 , 
        \test_module/add_46/n152 , \test_module/add_46/n154 , \test_module/add_46/n156 , 
        \test_module/add_46/n158 , \test_module/add_46/n160 , \test_module/add_46/n162 , 
        \test_module/add_46/n164 , \test_module/add_46/n166 , \test_module/add_46/n168 , 
        \test_module/add_46/n170 , \test_module/add_46/n172 , \test_module/add_46/n174 , 
        \test_module/add_46/n176 , \test_module/add_46/n178 , \test_module/add_46/n180 , 
        \test_module/add_46/n182 , \test_module/add_46/n184 , \test_module/add_46/n186 , 
        \test_module/add_46/n188 , \test_module/add_46/n190 , \test_module/add_46/n192 , 
        \test_module/add_46/n194 , \test_module/add_46/n196 , \test_module/add_46/n198 , 
        \test_module/add_46/n200 , \test_module/add_46/n202 , \test_module/add_46/n204 , 
        \test_module/add_46/n206 , \test_module/add_46/n208 , \test_module/add_46/n210 , 
        \test_module/add_46/n212 , \test_module/add_46/n214 , \test_module/add_46/n216 , 
        \test_module/add_46/n218 , \test_module/add_41/n182 , \test_module/add_46/n220 , 
        \test_module/add_46/n222 , \test_module/add_46/n224 , \test_module/add_46/n226 , 
        \test_module/add_46/n228 , \test_module/add_46/n230 , \test_module/add_46/n232 , 
        \test_module/add_46/n234 , \test_module/add_46/n236 , \test_module/add_46/n238 , 
        \test_module/add_46/n240 , \test_module/add_46/n242 , \test_module/add_46/n244 , 
        \test_module/add_46/n246 , \test_module/add_46/n248 , \test_module/add_46/n250 , 
        \test_module/add_46/n252 , \test_module/add_46/n254 , \test_module/add_46/n256 , 
        \test_module/add_46/n258 , \test_module/add_46/n260 , \test_module/add_46/n262 , 
        \test_module/add_46/n264 , \test_module/add_46/n266 , \test_module/add_46/n268 , 
        \test_module/add_46/n270 , \test_module/add_46/n272 , \test_module/add_46/n274 , 
        \test_module/add_46/n276 , \test_module/add_46/n278 , \test_module/add_46/n280 , 
        \test_module/add_46/n282 , \test_module/add_46/n284 , \test_module/add_46/n286 , 
        \test_module/add_46/n288 , \test_module/add_46/n290 , \test_module/add_46/n292 , 
        \test_module/add_46/n294 , \test_module/add_46/n296 , \test_module/add_46/n298 , 
        \test_module/add_46/n300 , \test_module/add_46/n302 , \test_module/add_46/n304 , 
        \test_module/add_46/n306 , \test_module/add_46/n308 , \test_module/add_46/n310 , 
        \test_module/add_46/n312 , \test_module/add_46/n314 , \test_module/add_46/n316 , 
        \test_module/add_46/n318 , \test_module/add_46/n320 , \test_module/add_46/n322 , 
        \test_module/add_46/n324 , \test_module/add_46/n326 , \test_module/add_46/n328 , 
        \test_module/add_46/n330 , \test_module/add_46/n332 , \test_module/add_46/n334 , 
        \test_module/add_46/n336 , \test_module/add_46/n338 , \test_module/add_46/n340 , 
        \test_module/add_46/n342 , \test_module/add_46/n344 , \test_module/add_46/n346 , 
        \test_module/add_46/n348 , \test_module/add_46/n350 , \test_module/add_46/n352 , 
        \test_module/add_46/n354 , \test_module/add_46/n356 , \test_module/add_46/n358 , 
        \test_module/add_46/n360 , \test_module/add_46/n362 , \test_module/add_46/n364 , 
        \test_module/add_46/n366 , \test_module/add_46/n368 , \test_module/add_46/n370 , 
        \test_module/add_46/n372 , \test_module/add_46/n374 , \test_module/add_46/n376 , 
        \test_module/add_46/n378 , \test_module/add_46/n380 , \test_module/add_46/n382 , 
        \test_module/add_46/n384 , \test_module/add_46/n386 , \test_module/add_46/n388 , 
        \test_module/add_46/n390 , \test_module/add_46/n392 , \test_module/add_46/n394 , 
        \test_module/add_46/n396 , \test_module/add_46/n398 , \test_module/add_46/n400 , 
        \test_module/add_46/n402 , \test_module/add_46/n404 , \test_module/add_46/n406 , 
        \test_module/add_46/n408 , \test_module/add_46/n410 , \test_module/add_46/n412 , 
        \test_module/add_46/n414 , \test_module/add_46/n416 , \test_module/add_46/n418 , 
        \test_module/add_46/n420 , \test_module/add_46/n422 , \test_module/add_46/n424 , 
        \test_module/add_46/n426 , \test_module/add_46/n428 , \test_module/add_46/n430 , 
        \test_module/add_46/n432 , \test_module/add_46/n434 , \test_module/add_46/n436 , 
        \test_module/add_46/n438 , \test_module/add_46/n440 , \test_module/add_46/n442 , 
        \test_module/add_46/n444 , \test_module/add_46/n446 , \test_module/add_46/n448 , 
        \test_module/add_46/n450 , \test_module/add_46/n452 , \test_module/add_46/n454 , 
        \test_module/add_46/n456 , \test_module/add_46/n458 , \test_module/add_46/n460 , 
        \test_module/add_46/n462 , \test_module/add_46/n464 , \test_module/add_46/n466 , 
        \test_module/add_46/n468 , \test_module/add_46/n470 , \test_module/add_46/n472 , 
        \test_module/add_46/n474 , \test_module/add_46/n476 , \test_module/add_46/n478 , 
        \test_module/add_46/n480 , \test_module/add_46/n482 , \test_module/add_46/n484 , 
        \test_module/add_46/n486 , \test_module/add_46/n488 , \test_module/add_46/n490 , 
        \test_module/add_46/n492 , \test_module/add_46/n494 , \test_module/add_46/n496 , 
        \test_module/add_46/n498 , \test_module/add_46/n500 , \test_module/add_46/n502 , 
        \test_module/add_46/n504 , \test_module/add_46/n506 , \test_module/add_46/n508 , 
        \debug_inst/vio0/vio_core_inst/add_772/n4 , \debug_inst/vio0/vio_core_inst/add_772/n6 , 
        \debug_inst/vio0/vio_core_inst/add_772/n8 , \debug_inst/vio0/vio_core_inst/add_33/n6 , 
        \debug_inst/vio0/vio_core_inst/add_33/n8 , \debug_inst/vio0/vio_core_inst/add_33/n10 ;
    wire [3:0]\debug_inst/vio0/vio_core_inst/opcode ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1188)
    wire [31:0]\debug_inst/vio0/vio_core_inst/address_counter ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1189)
    
    wire \test_module/add_41/n100 , \test_module/add_41/n98 , \test_module/add_41/n96 , 
        \test_module/add_41/n94 , \test_module/add_41/n92 , \test_module/add_41/n90 , 
        \test_module/add_41/n88 , \test_module/add_41/n86 , \test_module/add_41/n84 , 
        \test_module/add_41/n82 , \debug_inst/vio0/vio_core_inst/commit_sync1 , 
        \debug_inst/vio0/vio_core_inst/commit_sync2 , i_reg_rstn;
    wire [0:0]\debug_inst/vio0/vio_core_inst/probe_out_sync ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1256)
    
    wire \test_module/add_41/n80 ;
    wire [3:0]\debug_inst/vio0/vio_core_inst/internal_register_select ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1187)
    
    wire \test_module/add_41/n78 , \test_module/add_41/n174 , \test_module/add_41/n76 , 
        \test_module/add_41/n74 , \test_module/add_41/n72 , \test_module/add_41/n70 , 
        \test_module/add_41/n68 , \test_module/add_41/n66 , \test_module/add_41/n64 , 
        \test_module/add_41/n62 , \test_module/add_41/n60 , \test_module/add_41/n58 , 
        \test_module/add_41/n56 , \test_module/add_41/n54 , \test_module/add_41/n52 , 
        \test_module/add_41/n50 , \test_module/add_41/n48 , \test_module/add_41/n46 , 
        \test_module/add_41/n44 , \test_module/add_41/n42 , \test_module/add_41/n40 , 
        \test_module/add_41/n38 , \test_module/add_41/n36 , \test_module/add_41/n34 , 
        \test_module/add_41/n32 , \test_module/add_41/n30 , \test_module/add_41/n28 , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clkb ;
    wire [511:0]\debug_inst/vio0/vio_core_inst/probe_in_sync ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1253)
    
    wire \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clkb , 
        \test_module/add_41/n26 , \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clka , 
        \test_module/add_41/n24 , \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clka , 
        \test_module/add_41/n22 , \test_module/add_41/n20 , \test_module/add_41/n18 , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clkb , 
        \test_module/add_41/n16 , \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clka , 
        \test_module/add_41/n14 , \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clka , 
        \test_module/add_41/n12 , \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clka , 
        \test_module/add_41/n10 , \test_module/add_41/n8 , \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clkb , 
        \test_module/add_41/n6 , \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clka , 
        \test_module/add_41/n4 , \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clka ;
    wire [20:0]\test_module/n9 ;
    
    wire \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clkb , 
        \test_module/add_39/n24 , \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clka , 
        \test_module/add_39/n22 , \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clka , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clkb , 
        \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clka , 
        \test_module/add_39/n20 , \test_module/add_39/n18 , \test_module/add_39/n16 , 
        \test_module/add_39/n14 , \test_module/add_39/n12 , \test_module/add_39/n10 , 
        \test_module/add_39/n8 , \test_module/add_39/n6 , \test_module/add_39/n4 ;
    wire [3:0]\debug_inst/debug_hub_inst/module_id_reg ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(410)
    
    wire \debug_inst/edb_soft_reset , \test_module/add_41/n188 , \test_module/add_41/n186 , 
        \test_module/add_39/n2 ;
    wire [81:0]\debug_inst/edb_user_dr ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(34)
    wire [20:0]\test_module/n569 ;
    
    wire ceg_net2, \~test_module/equal_21/n41 ;
    wire [20:0]\test_module/n1692 ;
    
    wire ceg_net5, \~test_module/equal_8/n41 , \debug_inst/vio0/vio_core_inst/n251 , 
        \clk_1~O ;
    wire [5:0]\debug_inst/vio0/vio_core_inst/n422 ;
    
    wire ceg_net8, \debug_inst/vio0/vio_core_inst/addr_ct_en ;
    wire [15:0]\debug_inst/vio0/vio_core_inst/data_to_word_counter ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1239)
    
    wire \debug_inst/vio0/vio_core_inst/word_ct_en ;
    wire [15:0]\debug_inst/vio0/vio_core_inst/n546 ;
    
    wire ceg_net11;
    wire [3:0]\debug_inst/vio0/vio_core_inst/module_next_state ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1246)
    wire [15:0]\debug_inst/vio0/vio_core_inst/probe_in_mux_out ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1824)
    
    wire \debug_inst/vio0/vio_core_inst/n2907 ;
    wire [31:0]\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 ;
    
    wire ceg_net16, \debug_inst/vio0/vio_core_inst/op_reg_en ;
    wire [31:0]\debug_inst/vio0/vio_core_inst/data_to_addr_counter ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1236)
    
    wire \debug_inst/vio0/vio_core_inst/n2952 , \debug_inst/vio0/vio_core_inst/regsel_ld_en , 
        \debug_inst/debug_hub_inst/n267 , \debug_inst/debug_hub_inst/n265 , 
        \clk_0~O , \debug_inst/debug_hub_inst/n96 , \bscan_TCK~O , n4093, 
        n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, 
        n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, 
        n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, 
        n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, 
        n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, 
        n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, 
        n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, 
        n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, 
        n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, 
        n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, 
        n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, 
        n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, 
        n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, 
        n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, 
        n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, 
        n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, 
        n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, 
        n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, 
        n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, 
        n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, 
        n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, 
        n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, 
        n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, 
        n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, 
        n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, 
        n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, 
        n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, 
        n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, 
        n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, 
        n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, 
        n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, 
        n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, 
        n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, 
        n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, 
        n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, 
        n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, 
        n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, 
        n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, 
        n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, 
        n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, 
        n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, 
        n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, 
        n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, 
        n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, 
        n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, 
        n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, 
        n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, 
        n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, 
        n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, 
        n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, 
        n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, 
        n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, 
        n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, 
        n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, 
        n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, 
        n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, 
        n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, 
        n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, 
        n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, 
        n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, 
        n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, 
        n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, 
        n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, 
        n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, 
        n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, 
        n4614;
    
    EFX_LUT4 LUT__10217 (.I0(\debug_inst/vio0/vio_core_inst/crc_data_out [24]), 
            .I1(\debug_inst/edb_user_dr [74]), .I2(\debug_inst/edb_user_dr [54]), 
            .I3(\debug_inst/vio0/vio_core_inst/crc_data_out [4]), .O(n4093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__10217.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__10218 (.I0(\debug_inst/vio0/vio_core_inst/crc_data_out [28]), 
            .I1(\debug_inst/edb_user_dr [78]), .I2(\debug_inst/edb_user_dr [70]), 
            .I3(\debug_inst/vio0/vio_core_inst/crc_data_out [20]), .O(n4094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__10218.LUTMASK = 16'h9009;
    EFX_FF \test_module/delay_1[0]~FF  (.D(\test_module/n569 [0]), .CE(ceg_net2), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(\test_module/delay_1 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \test_module/delay_1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_1[0]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_1[0]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_1[0]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_1[0]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_1[0]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[0]~FF  (.D(o_pllBr1_reg[0]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[0]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[0]~FF .D_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_2[0]~FF  (.D(\test_module/n1692 [0]), .CE(ceg_net5), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(\test_module/delay_2 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \test_module/delay_2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_2[0]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_2[0]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_2[0]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_2[0]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_2[0]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[1]~FF  (.D(\test_module/n33 [1]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[1]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[0]~FF  (.D(o_pllBr0_reg[0]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[0]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[0]~FF .D_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_1[1]~FF  (.D(\test_module/n569 [1]), .CE(ceg_net2), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(\test_module/delay_1 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \test_module/delay_1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_1[1]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_1[1]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_1[1]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_1[1]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_1[1]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_1[2]~FF  (.D(\test_module/n569 [2]), .CE(ceg_net2), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(\test_module/delay_1 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \test_module/delay_1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_1[2]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_1[2]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_1[2]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_1[2]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_1[2]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_1[3]~FF  (.D(\test_module/n569 [3]), .CE(ceg_net2), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(\test_module/delay_1 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \test_module/delay_1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_1[3]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_1[3]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_1[3]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_1[3]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_1[3]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_1[4]~FF  (.D(\test_module/n569 [4]), .CE(ceg_net2), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(\test_module/delay_1 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \test_module/delay_1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_1[4]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_1[4]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_1[4]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_1[4]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_1[4]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_1[5]~FF  (.D(\test_module/n569 [5]), .CE(ceg_net2), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(\test_module/delay_1 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \test_module/delay_1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_1[5]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_1[5]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_1[5]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_1[5]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_1[5]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_1[6]~FF  (.D(\test_module/n569 [6]), .CE(ceg_net2), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(\test_module/delay_1 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \test_module/delay_1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_1[6]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_1[6]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_1[6]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_1[6]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_1[6]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_1[7]~FF  (.D(\test_module/n569 [7]), .CE(ceg_net2), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(\test_module/delay_1 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \test_module/delay_1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_1[7]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_1[7]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_1[7]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_1[7]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_1[7]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_1[8]~FF  (.D(\test_module/n569 [8]), .CE(ceg_net2), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(\test_module/delay_1 [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \test_module/delay_1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_1[8]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_1[8]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_1[8]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_1[8]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_1[8]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_1[9]~FF  (.D(\test_module/n569 [9]), .CE(ceg_net2), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(\test_module/delay_1 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \test_module/delay_1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_1[9]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_1[9]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_1[9]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_1[9]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_1[9]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_1[10]~FF  (.D(\test_module/n569 [10]), .CE(ceg_net2), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(\test_module/delay_1 [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \test_module/delay_1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_1[10]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_1[10]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_1[10]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_1[10]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_1[10]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_1[11]~FF  (.D(\test_module/n569 [11]), .CE(ceg_net2), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(\test_module/delay_1 [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \test_module/delay_1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_1[11]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_1[11]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_1[11]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_1[11]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_1[11]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_1[12]~FF  (.D(\test_module/n569 [12]), .CE(ceg_net2), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(\test_module/delay_1 [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \test_module/delay_1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_1[12]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_1[12]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_1[12]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_1[12]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_1[12]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_1[13]~FF  (.D(\test_module/n569 [13]), .CE(ceg_net2), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(\test_module/delay_1 [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \test_module/delay_1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_1[13]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_1[13]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_1[13]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_1[13]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_1[13]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[1]~FF  (.D(\test_module/n1156 [1]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[1]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[2]~FF  (.D(\test_module/n1156 [2]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[2]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[3]~FF  (.D(\test_module/n1156 [3]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[3]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[4]~FF  (.D(\test_module/n1156 [4]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[4]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[4]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[5]~FF  (.D(\test_module/n1156 [5]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[5]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[5]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[5]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[6]~FF  (.D(\test_module/n1156 [6]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[6]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[6]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[6]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[7]~FF  (.D(\test_module/n1156 [7]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[7]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[7]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[7]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[8]~FF  (.D(\test_module/n1156 [8]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[8]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[8]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[8]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[8]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[8]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[8]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[9]~FF  (.D(\test_module/n1156 [9]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[9]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[9]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[9]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[9]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[9]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[9]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[10]~FF  (.D(\test_module/n1156 [10]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[10]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[10]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[10]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[10]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[10]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[10]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[11]~FF  (.D(\test_module/n1156 [11]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[11]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[11]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[11]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[11]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[11]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[11]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[12]~FF  (.D(\test_module/n1156 [12]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[12]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[12]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[12]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[12]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[12]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[12]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[13]~FF  (.D(\test_module/n1156 [13]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[13]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[13]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[13]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[13]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[13]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[13]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[14]~FF  (.D(\test_module/n1156 [14]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[14]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[14]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[14]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[14]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[14]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[14]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[15]~FF  (.D(\test_module/n1156 [15]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[15]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[15]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[16]~FF  (.D(\test_module/n1156 [16]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[16]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[16]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[17]~FF  (.D(\test_module/n1156 [17]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[17]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[17]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[18]~FF  (.D(\test_module/n1156 [18]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[18]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[18]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[19]~FF  (.D(\test_module/n1156 [19]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[19]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[19]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[20]~FF  (.D(\test_module/n1156 [20]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[20]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[20]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[21]~FF  (.D(\test_module/n1156 [21]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[21]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[21]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[22]~FF  (.D(\test_module/n1156 [22]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[22]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[22]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[23]~FF  (.D(\test_module/n1156 [23]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[23]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[23]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[24]~FF  (.D(\test_module/n1156 [24]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[24]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[24]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[25]~FF  (.D(\test_module/n1156 [25]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[25]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[25]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[25]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[25]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[25]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[25]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[26]~FF  (.D(\test_module/n1156 [26]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[26]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[26]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[26]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[26]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[26]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[26]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[27]~FF  (.D(\test_module/n1156 [27]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[27]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[27]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[27]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[27]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[27]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[27]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[28]~FF  (.D(\test_module/n1156 [28]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[28]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[28]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[28]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[28]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[28]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[28]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[29]~FF  (.D(\test_module/n1156 [29]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[29]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[29]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[29]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[29]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[29]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[29]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[30]~FF  (.D(\test_module/n1156 [30]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[30]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[30]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[30]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[30]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[30]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[30]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[31]~FF  (.D(\test_module/n1156 [31]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[31]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[31]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[31]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[31]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[31]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[31]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[32]~FF  (.D(\test_module/n1156 [32]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[32]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[32]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[32]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[32]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[32]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[32]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[33]~FF  (.D(\test_module/n1156 [33]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[33]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[33]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[33]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[33]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[33]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[33]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[34]~FF  (.D(\test_module/n1156 [34]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[34]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[34]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[34]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[34]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[34]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[34]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[35]~FF  (.D(\test_module/n1156 [35]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[35]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[35]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[35]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[35]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[35]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[35]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[36]~FF  (.D(\test_module/n1156 [36]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[36]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[36]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[36]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[36]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[36]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[36]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[37]~FF  (.D(\test_module/n1156 [37]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[37]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[37]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[37]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[37]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[37]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[37]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[38]~FF  (.D(\test_module/n1156 [38]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[38]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[38]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[38]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[38]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[38]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[38]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[39]~FF  (.D(\test_module/n1156 [39]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[39]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[39]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[39]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[39]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[39]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[39]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[40]~FF  (.D(\test_module/n1156 [40]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[40]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[40]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[40]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[40]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[40]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[40]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[41]~FF  (.D(\test_module/n1156 [41]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[41]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[41]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[41]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[41]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[41]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[41]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[42]~FF  (.D(\test_module/n1156 [42]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[42]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[42]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[42]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[42]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[42]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[42]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[43]~FF  (.D(\test_module/n1156 [43]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[43]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[43]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[43]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[43]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[43]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[43]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[44]~FF  (.D(\test_module/n1156 [44]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[44]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[44]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[44]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[44]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[44]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[44]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[45]~FF  (.D(\test_module/n1156 [45]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[45]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[45]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[45]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[45]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[45]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[45]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[46]~FF  (.D(\test_module/n1156 [46]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[46]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[46]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[46]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[46]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[46]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[46]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[47]~FF  (.D(\test_module/n1156 [47]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[47]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[47]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[47]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[47]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[47]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[47]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[48]~FF  (.D(\test_module/n1156 [48]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[48]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[48]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[48]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[48]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[48]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[48]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[49]~FF  (.D(\test_module/n1156 [49]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[49]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[49]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[49]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[49]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[49]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[49]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[50]~FF  (.D(\test_module/n1156 [50]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[50]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[50]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[50]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[50]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[50]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[50]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[51]~FF  (.D(\test_module/n1156 [51]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[51]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[51]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[51]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[51]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[51]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[51]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[52]~FF  (.D(\test_module/n1156 [52]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[52]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[52]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[52]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[52]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[52]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[52]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[53]~FF  (.D(\test_module/n1156 [53]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[53]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[53]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[53]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[53]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[53]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[53]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[54]~FF  (.D(\test_module/n1156 [54]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[54]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[54]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[54]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[54]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[54]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[54]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[55]~FF  (.D(\test_module/n1156 [55]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[55]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[55]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[55]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[55]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[55]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[55]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[56]~FF  (.D(\test_module/n1156 [56]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[56]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[56]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[56]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[56]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[56]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[56]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[57]~FF  (.D(\test_module/n1156 [57]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[57]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[57]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[57]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[57]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[57]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[57]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[58]~FF  (.D(\test_module/n1156 [58]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[58]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[58]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[58]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[58]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[58]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[58]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[59]~FF  (.D(\test_module/n1156 [59]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[59]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[59]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[59]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[59]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[59]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[59]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[60]~FF  (.D(\test_module/n1156 [60]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[60])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[60]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[60]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[60]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[60]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[60]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[60]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[61]~FF  (.D(\test_module/n1156 [61]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[61])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[61]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[61]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[61]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[61]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[61]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[61]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[62]~FF  (.D(\test_module/n1156 [62]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[62])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[62]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[62]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[62]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[62]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[62]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[62]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[63]~FF  (.D(\test_module/n1156 [63]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[63]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[63]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[63]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[63]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[63]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[63]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[64]~FF  (.D(\test_module/n1156 [64]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[64])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[64]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[64]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[64]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[64]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[64]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[64]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[65]~FF  (.D(\test_module/n1156 [65]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[65])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[65]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[65]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[65]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[65]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[65]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[65]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[66]~FF  (.D(\test_module/n1156 [66]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[66])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[66]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[66]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[66]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[66]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[66]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[66]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[67]~FF  (.D(\test_module/n1156 [67]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[67])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[67]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[67]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[67]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[67]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[67]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[67]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[68]~FF  (.D(\test_module/n1156 [68]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[68])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[68]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[68]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[68]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[68]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[68]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[68]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[69]~FF  (.D(\test_module/n1156 [69]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[69])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[69]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[69]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[69]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[69]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[69]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[69]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[70]~FF  (.D(\test_module/n1156 [70]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[70])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[70]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[70]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[70]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[70]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[70]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[70]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[71]~FF  (.D(\test_module/n1156 [71]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[71])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[71]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[71]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[71]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[71]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[71]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[71]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[72]~FF  (.D(\test_module/n1156 [72]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[72])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[72]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[72]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[72]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[72]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[72]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[72]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[73]~FF  (.D(\test_module/n1156 [73]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[73])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[73]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[73]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[73]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[73]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[73]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[73]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[74]~FF  (.D(\test_module/n1156 [74]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[74])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[74]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[74]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[74]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[74]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[74]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[74]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[75]~FF  (.D(\test_module/n1156 [75]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[75])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[75]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[75]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[75]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[75]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[75]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[75]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[76]~FF  (.D(\test_module/n1156 [76]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[76])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[76]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[76]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[76]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[76]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[76]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[76]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[77]~FF  (.D(\test_module/n1156 [77]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[77])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[77]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[77]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[77]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[77]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[77]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[77]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[78]~FF  (.D(\test_module/n1156 [78]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[78])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[78]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[78]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[78]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[78]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[78]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[78]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[79]~FF  (.D(\test_module/n1156 [79]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[79])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[79]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[79]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[79]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[79]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[79]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[79]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[80]~FF  (.D(\test_module/n1156 [80]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[80])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[80]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[80]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[80]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[80]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[80]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[80]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[81]~FF  (.D(\test_module/n1156 [81]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[81])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[81]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[81]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[81]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[81]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[81]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[81]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[82]~FF  (.D(\test_module/n1156 [82]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[82])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[82]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[82]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[82]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[82]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[82]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[82]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[83]~FF  (.D(\test_module/n1156 [83]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[83])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[83]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[83]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[83]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[83]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[83]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[83]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[84]~FF  (.D(\test_module/n1156 [84]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[84])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[84]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[84]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[84]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[84]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[84]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[84]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[85]~FF  (.D(\test_module/n1156 [85]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[85])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[85]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[85]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[85]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[85]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[85]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[85]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[86]~FF  (.D(\test_module/n1156 [86]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[86])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[86]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[86]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[86]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[86]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[86]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[86]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[87]~FF  (.D(\test_module/n1156 [87]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[87])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[87]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[87]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[87]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[87]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[87]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[87]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[88]~FF  (.D(\test_module/n1156 [88]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[88])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[88]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[88]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[88]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[88]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[88]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[88]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[89]~FF  (.D(\test_module/n1156 [89]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[89])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[89]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[89]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[89]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[89]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[89]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[89]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[90]~FF  (.D(\test_module/n1156 [90]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[90])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[90]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[90]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[90]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[90]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[90]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[90]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[91]~FF  (.D(\test_module/n1156 [91]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[91])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[91]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[91]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[91]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[91]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[91]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[91]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[92]~FF  (.D(\test_module/n1156 [92]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[92])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[92]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[92]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[92]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[92]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[92]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[92]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[93]~FF  (.D(\test_module/n1156 [93]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[93])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[93]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[93]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[93]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[93]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[93]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[93]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[94]~FF  (.D(\test_module/n1156 [94]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[94])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[94]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[94]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[94]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[94]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[94]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[94]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[95]~FF  (.D(\test_module/n1156 [95]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[95])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[95]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[95]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[95]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[95]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[95]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[95]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[96]~FF  (.D(\test_module/n1156 [96]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[96])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[96]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[96]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[96]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[96]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[96]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[96]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[97]~FF  (.D(\test_module/n1156 [97]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[97])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[97]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[97]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[97]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[97]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[97]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[97]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[98]~FF  (.D(\test_module/n1156 [98]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[98])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[98]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[98]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[98]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[98]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[98]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[98]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[99]~FF  (.D(\test_module/n1156 [99]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[99])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[99]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[99]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[99]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[99]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[99]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[99]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[100]~FF  (.D(\test_module/n1156 [100]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[100])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[100]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[100]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[100]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[100]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[100]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[100]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[101]~FF  (.D(\test_module/n1156 [101]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[101])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[101]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[101]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[101]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[101]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[101]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[101]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[102]~FF  (.D(\test_module/n1156 [102]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[102])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[102]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[102]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[102]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[102]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[102]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[102]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[103]~FF  (.D(\test_module/n1156 [103]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[103])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[103]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[103]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[103]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[103]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[103]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[103]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[104]~FF  (.D(\test_module/n1156 [104]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[104])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[104]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[104]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[104]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[104]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[104]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[104]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[105]~FF  (.D(\test_module/n1156 [105]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[105])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[105]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[105]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[105]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[105]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[105]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[105]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[106]~FF  (.D(\test_module/n1156 [106]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[106])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[106]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[106]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[106]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[106]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[106]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[106]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[107]~FF  (.D(\test_module/n1156 [107]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[107])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[107]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[107]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[107]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[107]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[107]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[107]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[108]~FF  (.D(\test_module/n1156 [108]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[108])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[108]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[108]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[108]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[108]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[108]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[108]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[109]~FF  (.D(\test_module/n1156 [109]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[109])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[109]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[109]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[109]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[109]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[109]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[109]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[110]~FF  (.D(\test_module/n1156 [110]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[110])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[110]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[110]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[110]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[110]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[110]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[110]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[111]~FF  (.D(\test_module/n1156 [111]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[111])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[111]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[111]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[111]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[111]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[111]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[111]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[112]~FF  (.D(\test_module/n1156 [112]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[112])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[112]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[112]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[112]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[112]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[112]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[112]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[113]~FF  (.D(\test_module/n1156 [113]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[113])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[113]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[113]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[113]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[113]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[113]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[113]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[114]~FF  (.D(\test_module/n1156 [114]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[114])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[114]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[114]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[114]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[114]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[114]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[114]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[115]~FF  (.D(\test_module/n1156 [115]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[115])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[115]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[115]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[115]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[115]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[115]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[115]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[116]~FF  (.D(\test_module/n1156 [116]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[116])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[116]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[116]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[116]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[116]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[116]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[116]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[117]~FF  (.D(\test_module/n1156 [117]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[117])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[117]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[117]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[117]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[117]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[117]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[117]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[118]~FF  (.D(\test_module/n1156 [118]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[118])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[118]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[118]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[118]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[118]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[118]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[118]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[119]~FF  (.D(\test_module/n1156 [119]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[119])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[119]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[119]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[119]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[119]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[119]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[119]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[120]~FF  (.D(\test_module/n1156 [120]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[120])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[120]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[120]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[120]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[120]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[120]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[120]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[120]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[121]~FF  (.D(\test_module/n1156 [121]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[121])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[121]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[121]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[121]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[121]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[121]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[121]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[121]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[122]~FF  (.D(\test_module/n1156 [122]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[122])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[122]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[122]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[122]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[122]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[122]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[122]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[122]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[123]~FF  (.D(\test_module/n1156 [123]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[123])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[123]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[123]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[123]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[123]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[123]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[123]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[123]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[124]~FF  (.D(\test_module/n1156 [124]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[124])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[124]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[124]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[124]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[124]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[124]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[124]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[124]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[125]~FF  (.D(\test_module/n1156 [125]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[125])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[125]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[125]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[125]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[125]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[125]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[125]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[125]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[126]~FF  (.D(\test_module/n1156 [126]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[126])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[126]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[126]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[126]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[126]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[126]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[126]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[126]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[127]~FF  (.D(\test_module/n1156 [127]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[127])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[127]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[127]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[127]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[127]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[127]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[127]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[127]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[128]~FF  (.D(\test_module/n1156 [128]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[128])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[128]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[128]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[128]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[128]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[128]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[128]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[128]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[129]~FF  (.D(\test_module/n1156 [129]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[129])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[129]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[129]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[129]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[129]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[129]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[129]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[129]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[130]~FF  (.D(\test_module/n1156 [130]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[130])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[130]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[130]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[130]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[130]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[130]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[130]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[130]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[131]~FF  (.D(\test_module/n1156 [131]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[131])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[131]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[131]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[131]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[131]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[131]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[131]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[131]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[132]~FF  (.D(\test_module/n1156 [132]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[132])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[132]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[132]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[132]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[132]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[132]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[132]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[132]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[133]~FF  (.D(\test_module/n1156 [133]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[133])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[133]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[133]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[133]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[133]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[133]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[133]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[133]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[134]~FF  (.D(\test_module/n1156 [134]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[134])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[134]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[134]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[134]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[134]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[134]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[134]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[134]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[135]~FF  (.D(\test_module/n1156 [135]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[135])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[135]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[135]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[135]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[135]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[135]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[135]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[135]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[136]~FF  (.D(\test_module/n1156 [136]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[136])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[136]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[136]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[136]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[136]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[136]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[136]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[136]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[137]~FF  (.D(\test_module/n1156 [137]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[137])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[137]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[137]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[137]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[137]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[137]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[137]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[137]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[138]~FF  (.D(\test_module/n1156 [138]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[138])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[138]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[138]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[138]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[138]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[138]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[138]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[138]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[139]~FF  (.D(\test_module/n1156 [139]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[139])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[139]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[139]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[139]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[139]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[139]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[139]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[139]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[140]~FF  (.D(\test_module/n1156 [140]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[140])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[140]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[140]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[140]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[140]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[140]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[140]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[140]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[141]~FF  (.D(\test_module/n1156 [141]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[141])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[141]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[141]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[141]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[141]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[141]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[141]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[141]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[142]~FF  (.D(\test_module/n1156 [142]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[142])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[142]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[142]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[142]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[142]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[142]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[142]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[142]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[143]~FF  (.D(\test_module/n1156 [143]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[143])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[143]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[143]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[143]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[143]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[143]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[143]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[143]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[144]~FF  (.D(\test_module/n1156 [144]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[144])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[144]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[144]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[144]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[144]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[144]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[144]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[144]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[145]~FF  (.D(\test_module/n1156 [145]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[145])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[145]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[145]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[145]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[145]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[145]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[145]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[145]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[146]~FF  (.D(\test_module/n1156 [146]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[146])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[146]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[146]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[146]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[146]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[146]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[146]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[146]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[147]~FF  (.D(\test_module/n1156 [147]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[147])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[147]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[147]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[147]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[147]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[147]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[147]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[147]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[148]~FF  (.D(\test_module/n1156 [148]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[148])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[148]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[148]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[148]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[148]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[148]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[148]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[148]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[149]~FF  (.D(\test_module/n1156 [149]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[149])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[149]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[149]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[149]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[149]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[149]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[149]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[149]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[150]~FF  (.D(\test_module/n1156 [150]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[150])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[150]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[150]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[150]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[150]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[150]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[150]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[150]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[151]~FF  (.D(\test_module/n1156 [151]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[151])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[151]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[151]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[151]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[151]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[151]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[151]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[151]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[152]~FF  (.D(\test_module/n1156 [152]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[152])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[152]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[152]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[152]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[152]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[152]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[152]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[152]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[153]~FF  (.D(\test_module/n1156 [153]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[153])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[153]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[153]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[153]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[153]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[153]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[153]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[153]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[154]~FF  (.D(\test_module/n1156 [154]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[154])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[154]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[154]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[154]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[154]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[154]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[154]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[154]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[155]~FF  (.D(\test_module/n1156 [155]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[155])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[155]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[155]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[155]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[155]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[155]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[155]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[155]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[156]~FF  (.D(\test_module/n1156 [156]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[156])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[156]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[156]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[156]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[156]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[156]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[156]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[156]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[157]~FF  (.D(\test_module/n1156 [157]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[157])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[157]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[157]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[157]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[157]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[157]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[157]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[157]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[158]~FF  (.D(\test_module/n1156 [158]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[158])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[158]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[158]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[158]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[158]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[158]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[158]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[158]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[159]~FF  (.D(\test_module/n1156 [159]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[159])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[159]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[159]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[159]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[159]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[159]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[159]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[159]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[160]~FF  (.D(\test_module/n1156 [160]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[160])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[160]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[160]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[160]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[160]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[160]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[160]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[160]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[161]~FF  (.D(\test_module/n1156 [161]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[161])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[161]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[161]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[161]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[161]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[161]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[161]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[161]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[162]~FF  (.D(\test_module/n1156 [162]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[162])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[162]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[162]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[162]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[162]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[162]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[162]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[162]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[163]~FF  (.D(\test_module/n1156 [163]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[163])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[163]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[163]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[163]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[163]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[163]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[163]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[163]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[164]~FF  (.D(\test_module/n1156 [164]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[164])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[164]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[164]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[164]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[164]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[164]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[164]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[164]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[165]~FF  (.D(\test_module/n1156 [165]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[165])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[165]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[165]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[165]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[165]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[165]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[165]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[165]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[166]~FF  (.D(\test_module/n1156 [166]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[166])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[166]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[166]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[166]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[166]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[166]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[166]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[166]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[167]~FF  (.D(\test_module/n1156 [167]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[167])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[167]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[167]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[167]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[167]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[167]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[167]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[167]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[168]~FF  (.D(\test_module/n1156 [168]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[168])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[168]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[168]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[168]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[168]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[168]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[168]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[168]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[169]~FF  (.D(\test_module/n1156 [169]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[169])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[169]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[169]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[169]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[169]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[169]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[169]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[169]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[170]~FF  (.D(\test_module/n1156 [170]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[170])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[170]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[170]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[170]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[170]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[170]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[170]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[170]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[171]~FF  (.D(\test_module/n1156 [171]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[171])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[171]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[171]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[171]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[171]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[171]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[171]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[171]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[172]~FF  (.D(\test_module/n1156 [172]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[172])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[172]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[172]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[172]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[172]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[172]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[172]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[172]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[173]~FF  (.D(\test_module/n1156 [173]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[173])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[173]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[173]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[173]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[173]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[173]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[173]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[173]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[174]~FF  (.D(\test_module/n1156 [174]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[174])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[174]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[174]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[174]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[174]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[174]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[174]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[174]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[175]~FF  (.D(\test_module/n1156 [175]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[175])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[175]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[175]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[175]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[175]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[175]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[175]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[175]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[176]~FF  (.D(\test_module/n1156 [176]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[176])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[176]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[176]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[176]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[176]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[176]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[176]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[176]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[177]~FF  (.D(\test_module/n1156 [177]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[177])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[177]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[177]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[177]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[177]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[177]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[177]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[177]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[178]~FF  (.D(\test_module/n1156 [178]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[178])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[178]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[178]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[178]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[178]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[178]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[178]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[178]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[179]~FF  (.D(\test_module/n1156 [179]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[179])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[179]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[179]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[179]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[179]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[179]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[179]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[179]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[180]~FF  (.D(\test_module/n1156 [180]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[180])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[180]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[180]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[180]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[180]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[180]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[180]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[180]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[181]~FF  (.D(\test_module/n1156 [181]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[181])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[181]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[181]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[181]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[181]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[181]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[181]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[181]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[182]~FF  (.D(\test_module/n1156 [182]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[182])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[182]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[182]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[182]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[182]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[182]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[182]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[182]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[183]~FF  (.D(\test_module/n1156 [183]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[183])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[183]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[183]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[183]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[183]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[183]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[183]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[183]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[184]~FF  (.D(\test_module/n1156 [184]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[184])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[184]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[184]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[184]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[184]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[184]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[184]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[184]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[185]~FF  (.D(\test_module/n1156 [185]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[185])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[185]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[185]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[185]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[185]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[185]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[185]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[185]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[186]~FF  (.D(\test_module/n1156 [186]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[186])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[186]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[186]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[186]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[186]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[186]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[186]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[186]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[187]~FF  (.D(\test_module/n1156 [187]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[187])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[187]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[187]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[187]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[187]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[187]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[187]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[187]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[188]~FF  (.D(\test_module/n1156 [188]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[188])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[188]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[188]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[188]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[188]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[188]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[188]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[188]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[189]~FF  (.D(\test_module/n1156 [189]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[189])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[189]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[189]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[189]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[189]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[189]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[189]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[189]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[190]~FF  (.D(\test_module/n1156 [190]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[190])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[190]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[190]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[190]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[190]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[190]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[190]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[190]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[191]~FF  (.D(\test_module/n1156 [191]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[191])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[191]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[191]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[191]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[191]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[191]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[191]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[191]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[192]~FF  (.D(\test_module/n1156 [192]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[192])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[192]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[192]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[192]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[192]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[192]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[192]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[192]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[193]~FF  (.D(\test_module/n1156 [193]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[193])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[193]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[193]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[193]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[193]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[193]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[193]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[193]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[194]~FF  (.D(\test_module/n1156 [194]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[194])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[194]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[194]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[194]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[194]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[194]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[194]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[194]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[195]~FF  (.D(\test_module/n1156 [195]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[195])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[195]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[195]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[195]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[195]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[195]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[195]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[195]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[196]~FF  (.D(\test_module/n1156 [196]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[196])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[196]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[196]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[196]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[196]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[196]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[196]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[196]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[197]~FF  (.D(\test_module/n1156 [197]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[197])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[197]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[197]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[197]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[197]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[197]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[197]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[197]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[198]~FF  (.D(\test_module/n1156 [198]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[198])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[198]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[198]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[198]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[198]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[198]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[198]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[198]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[199]~FF  (.D(\test_module/n1156 [199]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[199])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[199]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[199]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[199]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[199]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[199]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[199]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[199]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[200]~FF  (.D(\test_module/n1156 [200]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[200])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[200]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[200]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[200]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[200]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[200]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[200]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[200]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[201]~FF  (.D(\test_module/n1156 [201]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[201])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[201]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[201]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[201]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[201]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[201]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[201]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[201]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[202]~FF  (.D(\test_module/n1156 [202]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[202])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[202]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[202]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[202]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[202]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[202]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[202]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[202]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[203]~FF  (.D(\test_module/n1156 [203]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[203])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[203]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[203]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[203]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[203]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[203]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[203]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[203]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[204]~FF  (.D(\test_module/n1156 [204]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[204])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[204]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[204]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[204]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[204]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[204]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[204]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[204]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[205]~FF  (.D(\test_module/n1156 [205]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[205])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[205]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[205]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[205]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[205]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[205]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[205]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[205]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[206]~FF  (.D(\test_module/n1156 [206]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[206])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[206]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[206]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[206]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[206]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[206]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[206]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[206]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[207]~FF  (.D(\test_module/n1156 [207]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[207])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[207]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[207]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[207]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[207]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[207]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[207]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[207]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[208]~FF  (.D(\test_module/n1156 [208]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[208])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[208]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[208]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[208]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[208]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[208]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[208]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[208]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[209]~FF  (.D(\test_module/n1156 [209]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[209])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[209]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[209]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[209]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[209]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[209]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[209]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[209]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[210]~FF  (.D(\test_module/n1156 [210]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[210])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[210]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[210]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[210]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[210]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[210]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[210]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[210]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[211]~FF  (.D(\test_module/n1156 [211]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[211])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[211]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[211]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[211]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[211]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[211]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[211]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[211]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[212]~FF  (.D(\test_module/n1156 [212]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[212])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[212]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[212]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[212]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[212]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[212]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[212]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[212]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[213]~FF  (.D(\test_module/n1156 [213]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[213])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[213]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[213]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[213]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[213]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[213]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[213]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[213]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[214]~FF  (.D(\test_module/n1156 [214]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[214])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[214]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[214]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[214]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[214]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[214]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[214]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[214]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[215]~FF  (.D(\test_module/n1156 [215]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[215])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[215]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[215]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[215]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[215]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[215]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[215]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[215]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[216]~FF  (.D(\test_module/n1156 [216]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[216])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[216]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[216]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[216]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[216]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[216]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[216]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[216]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[217]~FF  (.D(\test_module/n1156 [217]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[217])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[217]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[217]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[217]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[217]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[217]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[217]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[217]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[218]~FF  (.D(\test_module/n1156 [218]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[218])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[218]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[218]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[218]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[218]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[218]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[218]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[218]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[219]~FF  (.D(\test_module/n1156 [219]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[219])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[219]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[219]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[219]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[219]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[219]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[219]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[219]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[220]~FF  (.D(\test_module/n1156 [220]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[220])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[220]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[220]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[220]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[220]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[220]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[220]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[220]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[221]~FF  (.D(\test_module/n1156 [221]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[221])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[221]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[221]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[221]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[221]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[221]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[221]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[221]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[222]~FF  (.D(\test_module/n1156 [222]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[222])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[222]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[222]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[222]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[222]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[222]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[222]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[222]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[223]~FF  (.D(\test_module/n1156 [223]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[223])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[223]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[223]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[223]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[223]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[223]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[223]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[223]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[224]~FF  (.D(\test_module/n1156 [224]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[224])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[224]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[224]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[224]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[224]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[224]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[224]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[224]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[225]~FF  (.D(\test_module/n1156 [225]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[225])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[225]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[225]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[225]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[225]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[225]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[225]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[225]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[226]~FF  (.D(\test_module/n1156 [226]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[226])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[226]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[226]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[226]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[226]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[226]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[226]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[226]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[227]~FF  (.D(\test_module/n1156 [227]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[227])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[227]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[227]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[227]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[227]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[227]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[227]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[227]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[228]~FF  (.D(\test_module/n1156 [228]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[228])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[228]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[228]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[228]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[228]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[228]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[228]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[228]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[229]~FF  (.D(\test_module/n1156 [229]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[229])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[229]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[229]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[229]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[229]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[229]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[229]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[229]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[230]~FF  (.D(\test_module/n1156 [230]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[230])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[230]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[230]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[230]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[230]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[230]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[230]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[230]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[231]~FF  (.D(\test_module/n1156 [231]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[231])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[231]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[231]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[231]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[231]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[231]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[231]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[231]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[232]~FF  (.D(\test_module/n1156 [232]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[232])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[232]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[232]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[232]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[232]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[232]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[232]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[232]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[233]~FF  (.D(\test_module/n1156 [233]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[233])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[233]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[233]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[233]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[233]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[233]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[233]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[233]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[234]~FF  (.D(\test_module/n1156 [234]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[234])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[234]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[234]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[234]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[234]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[234]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[234]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[234]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[235]~FF  (.D(\test_module/n1156 [235]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[235])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[235]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[235]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[235]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[235]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[235]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[235]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[235]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[236]~FF  (.D(\test_module/n1156 [236]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[236])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[236]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[236]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[236]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[236]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[236]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[236]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[236]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[237]~FF  (.D(\test_module/n1156 [237]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[237])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[237]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[237]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[237]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[237]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[237]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[237]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[237]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[238]~FF  (.D(\test_module/n1156 [238]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[238])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[238]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[238]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[238]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[238]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[238]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[238]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[238]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[239]~FF  (.D(\test_module/n1156 [239]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[239])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[239]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[239]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[239]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[239]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[239]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[239]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[239]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[240]~FF  (.D(\test_module/n1156 [240]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[240])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[240]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[240]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[240]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[240]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[240]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[240]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[240]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[241]~FF  (.D(\test_module/n1156 [241]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[241])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[241]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[241]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[241]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[241]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[241]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[241]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[241]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[242]~FF  (.D(\test_module/n1156 [242]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[242])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[242]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[242]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[242]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[242]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[242]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[242]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[242]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[243]~FF  (.D(\test_module/n1156 [243]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[243])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[243]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[243]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[243]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[243]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[243]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[243]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[243]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[244]~FF  (.D(\test_module/n1156 [244]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[244])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[244]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[244]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[244]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[244]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[244]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[244]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[244]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[245]~FF  (.D(\test_module/n1156 [245]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[245])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[245]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[245]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[245]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[245]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[245]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[245]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[245]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[246]~FF  (.D(\test_module/n1156 [246]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[246])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[246]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[246]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[246]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[246]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[246]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[246]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[246]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[247]~FF  (.D(\test_module/n1156 [247]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[247])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[247]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[247]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[247]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[247]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[247]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[247]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[247]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[248]~FF  (.D(\test_module/n1156 [248]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[248])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[248]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[248]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[248]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[248]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[248]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[248]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[248]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[249]~FF  (.D(\test_module/n1156 [249]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[249])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[249]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[249]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[249]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[249]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[249]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[249]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[249]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[250]~FF  (.D(\test_module/n1156 [250]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[250])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[250]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[250]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[250]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[250]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[250]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[250]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[250]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[251]~FF  (.D(\test_module/n1156 [251]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[251])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[251]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[251]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[251]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[251]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[251]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[251]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[251]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[252]~FF  (.D(\test_module/n1156 [252]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[252])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[252]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[252]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[252]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[252]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[252]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[252]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[252]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[253]~FF  (.D(\test_module/n1156 [253]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[253])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[253]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[253]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[253]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[253]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[253]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[253]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[253]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[254]~FF  (.D(\test_module/n1156 [254]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[254])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[254]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[254]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[254]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[254]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[254]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[254]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[254]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr1_reg[255]~FF  (.D(\test_module/n1156 [255]), .CE(\~test_module/equal_21/n41 ), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(o_pllBr1_reg[255])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \o_pllBr1_reg[255]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[255]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[255]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr1_reg[255]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr1_reg[255]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr1_reg[255]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr1_reg[255]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_2[1]~FF  (.D(\test_module/n1692 [1]), .CE(ceg_net5), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(\test_module/delay_2 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \test_module/delay_2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_2[1]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_2[1]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_2[1]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_2[1]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_2[1]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_2[2]~FF  (.D(\test_module/n1692 [2]), .CE(ceg_net5), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(\test_module/delay_2 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \test_module/delay_2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_2[2]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_2[2]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_2[2]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_2[2]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_2[2]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_2[3]~FF  (.D(\test_module/n1692 [3]), .CE(ceg_net5), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(\test_module/delay_2 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \test_module/delay_2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_2[3]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_2[3]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_2[3]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_2[3]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_2[3]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_2[4]~FF  (.D(\test_module/n1692 [4]), .CE(ceg_net5), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(\test_module/delay_2 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \test_module/delay_2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_2[4]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_2[4]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_2[4]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_2[4]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_2[4]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_2[5]~FF  (.D(\test_module/n1692 [5]), .CE(ceg_net5), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(\test_module/delay_2 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \test_module/delay_2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_2[5]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_2[5]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_2[5]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_2[5]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_2[5]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_2[6]~FF  (.D(\test_module/n1692 [6]), .CE(ceg_net5), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(\test_module/delay_2 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \test_module/delay_2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_2[6]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_2[6]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_2[6]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_2[6]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_2[6]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_2[7]~FF  (.D(\test_module/n1692 [7]), .CE(ceg_net5), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(\test_module/delay_2 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \test_module/delay_2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_2[7]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_2[7]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_2[7]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_2[7]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_2[7]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_2[8]~FF  (.D(\test_module/n1692 [8]), .CE(ceg_net5), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(\test_module/delay_2 [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \test_module/delay_2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_2[8]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_2[8]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_2[8]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_2[8]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_2[8]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_2[9]~FF  (.D(\test_module/n1692 [9]), .CE(ceg_net5), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(\test_module/delay_2 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \test_module/delay_2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_2[9]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_2[9]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_2[9]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_2[9]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_2[9]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_2[10]~FF  (.D(\test_module/n1692 [10]), .CE(ceg_net5), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(\test_module/delay_2 [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \test_module/delay_2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_2[10]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_2[10]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_2[10]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_2[10]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_2[10]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_2[11]~FF  (.D(\test_module/n1692 [11]), .CE(ceg_net5), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(\test_module/delay_2 [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \test_module/delay_2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_2[11]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_2[11]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_2[11]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_2[11]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_2[11]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_2[12]~FF  (.D(\test_module/n1692 [12]), .CE(ceg_net5), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(\test_module/delay_2 [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \test_module/delay_2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_2[12]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_2[12]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_2[12]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_2[12]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_2[12]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \test_module/delay_2[13]~FF  (.D(\test_module/n1692 [13]), .CE(ceg_net5), 
           .CLK(\clk_1~O ), .SR(i_reg_rstn), .Q(\test_module/delay_2 [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(39)
    defparam \test_module/delay_2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \test_module/delay_2[13]~FF .CE_POLARITY = 1'b0;
    defparam \test_module/delay_2[13]~FF .SR_POLARITY = 1'b0;
    defparam \test_module/delay_2[13]~FF .D_POLARITY = 1'b1;
    defparam \test_module/delay_2[13]~FF .SR_SYNC = 1'b0;
    defparam \test_module/delay_2[13]~FF .SR_VALUE = 1'b0;
    defparam \test_module/delay_2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[2]~FF  (.D(\test_module/n33 [2]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[2]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[3]~FF  (.D(\test_module/n33 [3]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[3]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[4]~FF  (.D(\test_module/n33 [4]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[4]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[4]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[5]~FF  (.D(\test_module/n33 [5]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[5]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[5]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[5]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[6]~FF  (.D(\test_module/n33 [6]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[6]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[6]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[6]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[7]~FF  (.D(\test_module/n33 [7]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[7]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[7]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[7]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[8]~FF  (.D(\test_module/n33 [8]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[8]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[8]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[8]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[8]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[8]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[8]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[9]~FF  (.D(\test_module/n33 [9]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[9]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[9]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[9]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[9]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[9]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[9]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[10]~FF  (.D(\test_module/n33 [10]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[10]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[10]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[10]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[10]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[10]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[10]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[11]~FF  (.D(\test_module/n33 [11]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[11]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[11]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[11]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[11]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[11]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[11]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[12]~FF  (.D(\test_module/n33 [12]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[12]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[12]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[12]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[12]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[12]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[12]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[13]~FF  (.D(\test_module/n33 [13]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[13]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[13]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[13]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[13]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[13]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[13]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[14]~FF  (.D(\test_module/n33 [14]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[14]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[14]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[14]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[14]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[14]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[14]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[15]~FF  (.D(\test_module/n33 [15]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[15]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[15]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[16]~FF  (.D(\test_module/n33 [16]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[16]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[16]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[17]~FF  (.D(\test_module/n33 [17]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[17]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[17]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[18]~FF  (.D(\test_module/n33 [18]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[18]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[18]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[19]~FF  (.D(\test_module/n33 [19]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[19]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[19]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[20]~FF  (.D(\test_module/n33 [20]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[20]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[20]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[21]~FF  (.D(\test_module/n33 [21]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[21]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[21]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[22]~FF  (.D(\test_module/n33 [22]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[22]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[22]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[23]~FF  (.D(\test_module/n33 [23]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[23]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[23]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[24]~FF  (.D(\test_module/n33 [24]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[24]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[24]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[25]~FF  (.D(\test_module/n33 [25]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[25]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[25]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[25]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[25]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[25]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[25]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[26]~FF  (.D(\test_module/n33 [26]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[26]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[26]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[26]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[26]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[26]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[26]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[27]~FF  (.D(\test_module/n33 [27]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[27]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[27]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[27]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[27]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[27]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[27]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[28]~FF  (.D(\test_module/n33 [28]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[28]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[28]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[28]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[28]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[28]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[28]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[29]~FF  (.D(\test_module/n33 [29]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[29]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[29]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[29]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[29]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[29]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[29]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[30]~FF  (.D(\test_module/n33 [30]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[30]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[30]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[30]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[30]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[30]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[30]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[31]~FF  (.D(\test_module/n33 [31]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[31]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[31]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[31]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[31]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[31]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[31]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[32]~FF  (.D(\test_module/n33 [32]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[32]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[32]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[32]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[32]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[32]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[32]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[33]~FF  (.D(\test_module/n33 [33]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[33]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[33]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[33]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[33]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[33]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[33]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[34]~FF  (.D(\test_module/n33 [34]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[34]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[34]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[34]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[34]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[34]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[34]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[35]~FF  (.D(\test_module/n33 [35]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[35]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[35]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[35]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[35]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[35]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[35]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[36]~FF  (.D(\test_module/n33 [36]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[36]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[36]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[36]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[36]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[36]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[36]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[37]~FF  (.D(\test_module/n33 [37]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[37]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[37]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[37]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[37]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[37]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[37]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[38]~FF  (.D(\test_module/n33 [38]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[38]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[38]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[38]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[38]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[38]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[38]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[39]~FF  (.D(\test_module/n33 [39]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[39]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[39]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[39]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[39]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[39]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[39]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[40]~FF  (.D(\test_module/n33 [40]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[40]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[40]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[40]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[40]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[40]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[40]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[41]~FF  (.D(\test_module/n33 [41]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[41]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[41]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[41]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[41]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[41]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[41]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[42]~FF  (.D(\test_module/n33 [42]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[42]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[42]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[42]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[42]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[42]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[42]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[43]~FF  (.D(\test_module/n33 [43]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[43]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[43]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[43]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[43]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[43]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[43]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[44]~FF  (.D(\test_module/n33 [44]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[44]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[44]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[44]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[44]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[44]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[44]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[45]~FF  (.D(\test_module/n33 [45]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[45]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[45]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[45]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[45]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[45]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[45]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[46]~FF  (.D(\test_module/n33 [46]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[46]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[46]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[46]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[46]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[46]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[46]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[47]~FF  (.D(\test_module/n33 [47]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[47]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[47]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[47]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[47]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[47]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[47]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[48]~FF  (.D(\test_module/n33 [48]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[48]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[48]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[48]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[48]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[48]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[48]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[49]~FF  (.D(\test_module/n33 [49]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[49]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[49]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[49]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[49]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[49]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[49]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[50]~FF  (.D(\test_module/n33 [50]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[50]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[50]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[50]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[50]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[50]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[50]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[51]~FF  (.D(\test_module/n33 [51]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[51]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[51]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[51]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[51]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[51]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[51]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[52]~FF  (.D(\test_module/n33 [52]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[52]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[52]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[52]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[52]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[52]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[52]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[53]~FF  (.D(\test_module/n33 [53]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[53]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[53]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[53]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[53]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[53]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[53]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[54]~FF  (.D(\test_module/n33 [54]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[54]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[54]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[54]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[54]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[54]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[54]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[55]~FF  (.D(\test_module/n33 [55]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[55]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[55]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[55]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[55]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[55]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[55]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[56]~FF  (.D(\test_module/n33 [56]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[56]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[56]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[56]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[56]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[56]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[56]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[57]~FF  (.D(\test_module/n33 [57]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[57]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[57]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[57]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[57]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[57]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[57]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[58]~FF  (.D(\test_module/n33 [58]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[58]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[58]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[58]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[58]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[58]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[58]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[59]~FF  (.D(\test_module/n33 [59]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[59]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[59]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[59]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[59]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[59]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[59]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[60]~FF  (.D(\test_module/n33 [60]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[60])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[60]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[60]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[60]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[60]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[60]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[60]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[61]~FF  (.D(\test_module/n33 [61]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[61])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[61]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[61]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[61]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[61]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[61]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[61]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[62]~FF  (.D(\test_module/n33 [62]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[62])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[62]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[62]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[62]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[62]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[62]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[62]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[63]~FF  (.D(\test_module/n33 [63]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[63]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[63]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[63]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[63]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[63]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[63]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[64]~FF  (.D(\test_module/n33 [64]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[64])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[64]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[64]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[64]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[64]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[64]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[64]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[65]~FF  (.D(\test_module/n33 [65]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[65])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[65]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[65]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[65]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[65]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[65]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[65]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[66]~FF  (.D(\test_module/n33 [66]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[66])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[66]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[66]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[66]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[66]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[66]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[66]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[67]~FF  (.D(\test_module/n33 [67]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[67])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[67]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[67]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[67]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[67]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[67]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[67]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[68]~FF  (.D(\test_module/n33 [68]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[68])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[68]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[68]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[68]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[68]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[68]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[68]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[69]~FF  (.D(\test_module/n33 [69]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[69])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[69]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[69]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[69]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[69]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[69]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[69]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[70]~FF  (.D(\test_module/n33 [70]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[70])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[70]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[70]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[70]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[70]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[70]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[70]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[71]~FF  (.D(\test_module/n33 [71]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[71])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[71]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[71]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[71]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[71]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[71]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[71]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[72]~FF  (.D(\test_module/n33 [72]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[72])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[72]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[72]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[72]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[72]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[72]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[72]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[73]~FF  (.D(\test_module/n33 [73]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[73])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[73]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[73]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[73]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[73]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[73]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[73]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[74]~FF  (.D(\test_module/n33 [74]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[74])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[74]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[74]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[74]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[74]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[74]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[74]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[75]~FF  (.D(\test_module/n33 [75]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[75])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[75]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[75]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[75]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[75]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[75]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[75]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[76]~FF  (.D(\test_module/n33 [76]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[76])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[76]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[76]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[76]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[76]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[76]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[76]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[77]~FF  (.D(\test_module/n33 [77]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[77])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[77]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[77]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[77]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[77]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[77]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[77]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[78]~FF  (.D(\test_module/n33 [78]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[78])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[78]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[78]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[78]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[78]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[78]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[78]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[79]~FF  (.D(\test_module/n33 [79]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[79])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[79]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[79]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[79]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[79]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[79]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[79]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[80]~FF  (.D(\test_module/n33 [80]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[80])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[80]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[80]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[80]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[80]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[80]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[80]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[81]~FF  (.D(\test_module/n33 [81]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[81])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[81]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[81]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[81]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[81]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[81]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[81]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[82]~FF  (.D(\test_module/n33 [82]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[82])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[82]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[82]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[82]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[82]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[82]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[82]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[83]~FF  (.D(\test_module/n33 [83]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[83])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[83]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[83]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[83]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[83]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[83]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[83]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[84]~FF  (.D(\test_module/n33 [84]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[84])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[84]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[84]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[84]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[84]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[84]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[84]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[85]~FF  (.D(\test_module/n33 [85]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[85])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[85]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[85]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[85]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[85]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[85]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[85]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[86]~FF  (.D(\test_module/n33 [86]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[86])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[86]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[86]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[86]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[86]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[86]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[86]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[87]~FF  (.D(\test_module/n33 [87]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[87])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[87]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[87]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[87]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[87]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[87]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[87]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[88]~FF  (.D(\test_module/n33 [88]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[88])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[88]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[88]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[88]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[88]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[88]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[88]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[89]~FF  (.D(\test_module/n33 [89]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[89])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[89]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[89]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[89]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[89]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[89]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[89]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[90]~FF  (.D(\test_module/n33 [90]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[90])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[90]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[90]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[90]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[90]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[90]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[90]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[91]~FF  (.D(\test_module/n33 [91]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[91])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[91]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[91]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[91]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[91]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[91]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[91]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[92]~FF  (.D(\test_module/n33 [92]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[92])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[92]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[92]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[92]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[92]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[92]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[92]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[93]~FF  (.D(\test_module/n33 [93]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[93])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[93]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[93]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[93]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[93]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[93]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[93]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[94]~FF  (.D(\test_module/n33 [94]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[94])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[94]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[94]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[94]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[94]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[94]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[94]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[95]~FF  (.D(\test_module/n33 [95]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[95])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[95]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[95]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[95]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[95]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[95]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[95]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[96]~FF  (.D(\test_module/n33 [96]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[96])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[96]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[96]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[96]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[96]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[96]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[96]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[97]~FF  (.D(\test_module/n33 [97]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[97])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[97]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[97]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[97]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[97]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[97]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[97]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[98]~FF  (.D(\test_module/n33 [98]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[98])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[98]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[98]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[98]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[98]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[98]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[98]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[99]~FF  (.D(\test_module/n33 [99]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[99])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[99]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[99]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[99]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[99]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[99]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[99]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[100]~FF  (.D(\test_module/n33 [100]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[100])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[100]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[100]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[100]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[100]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[100]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[100]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[101]~FF  (.D(\test_module/n33 [101]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[101])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[101]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[101]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[101]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[101]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[101]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[101]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[102]~FF  (.D(\test_module/n33 [102]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[102])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[102]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[102]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[102]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[102]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[102]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[102]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[103]~FF  (.D(\test_module/n33 [103]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[103])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[103]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[103]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[103]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[103]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[103]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[103]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[104]~FF  (.D(\test_module/n33 [104]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[104])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[104]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[104]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[104]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[104]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[104]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[104]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[105]~FF  (.D(\test_module/n33 [105]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[105])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[105]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[105]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[105]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[105]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[105]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[105]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[106]~FF  (.D(\test_module/n33 [106]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[106])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[106]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[106]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[106]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[106]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[106]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[106]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[107]~FF  (.D(\test_module/n33 [107]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[107])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[107]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[107]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[107]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[107]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[107]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[107]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[108]~FF  (.D(\test_module/n33 [108]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[108])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[108]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[108]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[108]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[108]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[108]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[108]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[109]~FF  (.D(\test_module/n33 [109]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[109])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[109]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[109]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[109]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[109]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[109]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[109]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[110]~FF  (.D(\test_module/n33 [110]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[110])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[110]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[110]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[110]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[110]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[110]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[110]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[111]~FF  (.D(\test_module/n33 [111]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[111])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[111]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[111]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[111]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[111]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[111]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[111]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[112]~FF  (.D(\test_module/n33 [112]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[112])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[112]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[112]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[112]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[112]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[112]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[112]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[113]~FF  (.D(\test_module/n33 [113]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[113])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[113]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[113]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[113]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[113]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[113]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[113]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[114]~FF  (.D(\test_module/n33 [114]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[114])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[114]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[114]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[114]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[114]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[114]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[114]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[115]~FF  (.D(\test_module/n33 [115]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[115])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[115]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[115]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[115]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[115]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[115]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[115]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[116]~FF  (.D(\test_module/n33 [116]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[116])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[116]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[116]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[116]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[116]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[116]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[116]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[117]~FF  (.D(\test_module/n33 [117]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[117])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[117]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[117]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[117]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[117]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[117]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[117]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[118]~FF  (.D(\test_module/n33 [118]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[118])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[118]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[118]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[118]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[118]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[118]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[118]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[119]~FF  (.D(\test_module/n33 [119]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[119])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[119]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[119]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[119]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[119]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[119]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[119]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[120]~FF  (.D(\test_module/n33 [120]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[120])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[120]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[120]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[120]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[120]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[120]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[120]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[120]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[121]~FF  (.D(\test_module/n33 [121]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[121])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[121]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[121]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[121]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[121]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[121]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[121]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[121]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[122]~FF  (.D(\test_module/n33 [122]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[122])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[122]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[122]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[122]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[122]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[122]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[122]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[122]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[123]~FF  (.D(\test_module/n33 [123]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[123])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[123]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[123]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[123]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[123]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[123]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[123]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[123]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[124]~FF  (.D(\test_module/n33 [124]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[124])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[124]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[124]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[124]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[124]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[124]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[124]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[124]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[125]~FF  (.D(\test_module/n33 [125]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[125])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[125]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[125]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[125]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[125]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[125]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[125]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[125]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[126]~FF  (.D(\test_module/n33 [126]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[126])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[126]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[126]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[126]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[126]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[126]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[126]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[126]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[127]~FF  (.D(\test_module/n33 [127]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[127])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[127]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[127]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[127]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[127]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[127]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[127]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[127]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[128]~FF  (.D(\test_module/n33 [128]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[128])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[128]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[128]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[128]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[128]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[128]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[128]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[128]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[129]~FF  (.D(\test_module/n33 [129]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[129])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[129]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[129]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[129]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[129]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[129]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[129]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[129]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[130]~FF  (.D(\test_module/n33 [130]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[130])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[130]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[130]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[130]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[130]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[130]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[130]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[130]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[131]~FF  (.D(\test_module/n33 [131]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[131])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[131]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[131]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[131]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[131]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[131]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[131]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[131]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[132]~FF  (.D(\test_module/n33 [132]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[132])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[132]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[132]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[132]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[132]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[132]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[132]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[132]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[133]~FF  (.D(\test_module/n33 [133]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[133])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[133]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[133]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[133]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[133]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[133]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[133]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[133]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[134]~FF  (.D(\test_module/n33 [134]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[134])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[134]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[134]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[134]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[134]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[134]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[134]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[134]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[135]~FF  (.D(\test_module/n33 [135]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[135])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[135]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[135]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[135]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[135]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[135]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[135]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[135]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[136]~FF  (.D(\test_module/n33 [136]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[136])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[136]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[136]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[136]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[136]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[136]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[136]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[136]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[137]~FF  (.D(\test_module/n33 [137]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[137])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[137]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[137]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[137]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[137]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[137]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[137]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[137]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[138]~FF  (.D(\test_module/n33 [138]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[138])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[138]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[138]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[138]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[138]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[138]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[138]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[138]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[139]~FF  (.D(\test_module/n33 [139]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[139])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[139]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[139]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[139]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[139]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[139]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[139]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[139]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[140]~FF  (.D(\test_module/n33 [140]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[140])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[140]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[140]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[140]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[140]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[140]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[140]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[140]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[141]~FF  (.D(\test_module/n33 [141]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[141])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[141]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[141]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[141]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[141]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[141]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[141]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[141]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[142]~FF  (.D(\test_module/n33 [142]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[142])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[142]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[142]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[142]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[142]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[142]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[142]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[142]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[143]~FF  (.D(\test_module/n33 [143]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[143])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[143]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[143]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[143]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[143]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[143]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[143]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[143]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[144]~FF  (.D(\test_module/n33 [144]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[144])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[144]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[144]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[144]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[144]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[144]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[144]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[144]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[145]~FF  (.D(\test_module/n33 [145]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[145])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[145]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[145]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[145]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[145]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[145]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[145]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[145]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[146]~FF  (.D(\test_module/n33 [146]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[146])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[146]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[146]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[146]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[146]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[146]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[146]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[146]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[147]~FF  (.D(\test_module/n33 [147]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[147])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[147]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[147]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[147]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[147]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[147]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[147]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[147]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[148]~FF  (.D(\test_module/n33 [148]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[148])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[148]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[148]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[148]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[148]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[148]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[148]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[148]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[149]~FF  (.D(\test_module/n33 [149]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[149])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[149]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[149]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[149]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[149]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[149]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[149]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[149]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[150]~FF  (.D(\test_module/n33 [150]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[150])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[150]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[150]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[150]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[150]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[150]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[150]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[150]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[151]~FF  (.D(\test_module/n33 [151]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[151])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[151]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[151]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[151]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[151]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[151]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[151]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[151]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[152]~FF  (.D(\test_module/n33 [152]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[152])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[152]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[152]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[152]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[152]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[152]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[152]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[152]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[153]~FF  (.D(\test_module/n33 [153]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[153])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[153]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[153]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[153]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[153]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[153]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[153]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[153]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[154]~FF  (.D(\test_module/n33 [154]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[154])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[154]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[154]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[154]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[154]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[154]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[154]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[154]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[155]~FF  (.D(\test_module/n33 [155]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[155])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[155]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[155]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[155]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[155]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[155]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[155]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[155]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[156]~FF  (.D(\test_module/n33 [156]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[156])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[156]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[156]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[156]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[156]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[156]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[156]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[156]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[157]~FF  (.D(\test_module/n33 [157]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[157])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[157]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[157]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[157]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[157]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[157]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[157]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[157]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[158]~FF  (.D(\test_module/n33 [158]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[158])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[158]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[158]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[158]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[158]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[158]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[158]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[158]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[159]~FF  (.D(\test_module/n33 [159]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[159])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[159]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[159]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[159]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[159]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[159]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[159]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[159]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[160]~FF  (.D(\test_module/n33 [160]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[160])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[160]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[160]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[160]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[160]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[160]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[160]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[160]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[161]~FF  (.D(\test_module/n33 [161]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[161])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[161]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[161]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[161]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[161]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[161]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[161]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[161]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[162]~FF  (.D(\test_module/n33 [162]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[162])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[162]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[162]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[162]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[162]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[162]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[162]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[162]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[163]~FF  (.D(\test_module/n33 [163]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[163])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[163]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[163]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[163]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[163]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[163]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[163]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[163]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[164]~FF  (.D(\test_module/n33 [164]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[164])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[164]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[164]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[164]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[164]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[164]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[164]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[164]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[165]~FF  (.D(\test_module/n33 [165]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[165])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[165]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[165]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[165]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[165]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[165]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[165]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[165]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[166]~FF  (.D(\test_module/n33 [166]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[166])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[166]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[166]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[166]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[166]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[166]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[166]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[166]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[167]~FF  (.D(\test_module/n33 [167]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[167])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[167]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[167]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[167]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[167]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[167]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[167]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[167]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[168]~FF  (.D(\test_module/n33 [168]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[168])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[168]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[168]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[168]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[168]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[168]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[168]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[168]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[169]~FF  (.D(\test_module/n33 [169]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[169])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[169]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[169]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[169]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[169]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[169]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[169]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[169]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[170]~FF  (.D(\test_module/n33 [170]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[170])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[170]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[170]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[170]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[170]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[170]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[170]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[170]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[171]~FF  (.D(\test_module/n33 [171]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[171])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[171]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[171]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[171]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[171]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[171]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[171]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[171]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[172]~FF  (.D(\test_module/n33 [172]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[172])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[172]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[172]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[172]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[172]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[172]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[172]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[172]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[173]~FF  (.D(\test_module/n33 [173]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[173])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[173]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[173]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[173]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[173]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[173]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[173]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[173]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[174]~FF  (.D(\test_module/n33 [174]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[174])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[174]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[174]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[174]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[174]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[174]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[174]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[174]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[175]~FF  (.D(\test_module/n33 [175]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[175])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[175]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[175]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[175]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[175]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[175]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[175]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[175]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[176]~FF  (.D(\test_module/n33 [176]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[176])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[176]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[176]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[176]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[176]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[176]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[176]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[176]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[177]~FF  (.D(\test_module/n33 [177]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[177])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[177]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[177]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[177]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[177]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[177]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[177]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[177]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[178]~FF  (.D(\test_module/n33 [178]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[178])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[178]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[178]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[178]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[178]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[178]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[178]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[178]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[179]~FF  (.D(\test_module/n33 [179]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[179])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[179]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[179]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[179]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[179]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[179]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[179]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[179]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[180]~FF  (.D(\test_module/n33 [180]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[180])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[180]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[180]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[180]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[180]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[180]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[180]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[180]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[181]~FF  (.D(\test_module/n33 [181]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[181])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[181]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[181]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[181]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[181]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[181]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[181]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[181]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[182]~FF  (.D(\test_module/n33 [182]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[182])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[182]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[182]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[182]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[182]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[182]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[182]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[182]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[183]~FF  (.D(\test_module/n33 [183]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[183])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[183]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[183]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[183]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[183]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[183]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[183]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[183]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[184]~FF  (.D(\test_module/n33 [184]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[184])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[184]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[184]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[184]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[184]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[184]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[184]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[184]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[185]~FF  (.D(\test_module/n33 [185]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[185])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[185]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[185]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[185]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[185]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[185]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[185]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[185]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[186]~FF  (.D(\test_module/n33 [186]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[186])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[186]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[186]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[186]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[186]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[186]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[186]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[186]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[187]~FF  (.D(\test_module/n33 [187]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[187])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[187]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[187]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[187]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[187]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[187]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[187]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[187]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[188]~FF  (.D(\test_module/n33 [188]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[188])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[188]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[188]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[188]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[188]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[188]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[188]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[188]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[189]~FF  (.D(\test_module/n33 [189]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[189])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[189]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[189]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[189]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[189]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[189]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[189]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[189]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[190]~FF  (.D(\test_module/n33 [190]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[190])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[190]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[190]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[190]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[190]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[190]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[190]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[190]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[191]~FF  (.D(\test_module/n33 [191]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[191])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[191]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[191]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[191]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[191]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[191]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[191]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[191]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[192]~FF  (.D(\test_module/n33 [192]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[192])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[192]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[192]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[192]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[192]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[192]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[192]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[192]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[193]~FF  (.D(\test_module/n33 [193]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[193])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[193]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[193]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[193]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[193]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[193]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[193]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[193]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[194]~FF  (.D(\test_module/n33 [194]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[194])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[194]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[194]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[194]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[194]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[194]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[194]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[194]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[195]~FF  (.D(\test_module/n33 [195]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[195])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[195]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[195]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[195]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[195]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[195]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[195]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[195]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[196]~FF  (.D(\test_module/n33 [196]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[196])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[196]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[196]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[196]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[196]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[196]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[196]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[196]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[197]~FF  (.D(\test_module/n33 [197]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[197])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[197]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[197]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[197]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[197]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[197]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[197]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[197]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[198]~FF  (.D(\test_module/n33 [198]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[198])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[198]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[198]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[198]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[198]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[198]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[198]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[198]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[199]~FF  (.D(\test_module/n33 [199]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[199])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[199]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[199]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[199]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[199]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[199]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[199]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[199]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[200]~FF  (.D(\test_module/n33 [200]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[200])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[200]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[200]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[200]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[200]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[200]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[200]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[200]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[201]~FF  (.D(\test_module/n33 [201]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[201])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[201]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[201]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[201]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[201]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[201]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[201]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[201]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[202]~FF  (.D(\test_module/n33 [202]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[202])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[202]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[202]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[202]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[202]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[202]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[202]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[202]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[203]~FF  (.D(\test_module/n33 [203]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[203])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[203]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[203]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[203]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[203]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[203]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[203]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[203]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[204]~FF  (.D(\test_module/n33 [204]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[204])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[204]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[204]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[204]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[204]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[204]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[204]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[204]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[205]~FF  (.D(\test_module/n33 [205]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[205])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[205]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[205]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[205]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[205]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[205]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[205]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[205]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[206]~FF  (.D(\test_module/n33 [206]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[206])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[206]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[206]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[206]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[206]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[206]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[206]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[206]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[207]~FF  (.D(\test_module/n33 [207]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[207])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[207]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[207]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[207]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[207]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[207]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[207]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[207]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[208]~FF  (.D(\test_module/n33 [208]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[208])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[208]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[208]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[208]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[208]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[208]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[208]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[208]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[209]~FF  (.D(\test_module/n33 [209]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[209])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[209]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[209]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[209]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[209]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[209]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[209]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[209]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[210]~FF  (.D(\test_module/n33 [210]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[210])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[210]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[210]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[210]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[210]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[210]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[210]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[210]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[211]~FF  (.D(\test_module/n33 [211]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[211])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[211]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[211]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[211]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[211]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[211]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[211]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[211]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[212]~FF  (.D(\test_module/n33 [212]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[212])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[212]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[212]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[212]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[212]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[212]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[212]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[212]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[213]~FF  (.D(\test_module/n33 [213]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[213])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[213]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[213]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[213]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[213]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[213]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[213]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[213]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[214]~FF  (.D(\test_module/n33 [214]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[214])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[214]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[214]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[214]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[214]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[214]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[214]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[214]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[215]~FF  (.D(\test_module/n33 [215]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[215])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[215]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[215]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[215]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[215]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[215]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[215]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[215]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[216]~FF  (.D(\test_module/n33 [216]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[216])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[216]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[216]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[216]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[216]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[216]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[216]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[216]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[217]~FF  (.D(\test_module/n33 [217]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[217])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[217]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[217]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[217]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[217]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[217]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[217]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[217]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[218]~FF  (.D(\test_module/n33 [218]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[218])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[218]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[218]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[218]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[218]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[218]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[218]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[218]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[219]~FF  (.D(\test_module/n33 [219]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[219])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[219]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[219]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[219]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[219]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[219]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[219]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[219]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[220]~FF  (.D(\test_module/n33 [220]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[220])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[220]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[220]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[220]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[220]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[220]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[220]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[220]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[221]~FF  (.D(\test_module/n33 [221]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[221])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[221]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[221]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[221]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[221]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[221]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[221]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[221]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[222]~FF  (.D(\test_module/n33 [222]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[222])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[222]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[222]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[222]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[222]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[222]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[222]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[222]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[223]~FF  (.D(\test_module/n33 [223]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[223])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[223]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[223]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[223]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[223]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[223]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[223]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[223]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[224]~FF  (.D(\test_module/n33 [224]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[224])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[224]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[224]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[224]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[224]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[224]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[224]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[224]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[225]~FF  (.D(\test_module/n33 [225]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[225])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[225]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[225]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[225]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[225]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[225]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[225]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[225]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[226]~FF  (.D(\test_module/n33 [226]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[226])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[226]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[226]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[226]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[226]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[226]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[226]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[226]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[227]~FF  (.D(\test_module/n33 [227]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[227])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[227]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[227]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[227]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[227]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[227]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[227]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[227]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[228]~FF  (.D(\test_module/n33 [228]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[228])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[228]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[228]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[228]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[228]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[228]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[228]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[228]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[229]~FF  (.D(\test_module/n33 [229]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[229])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[229]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[229]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[229]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[229]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[229]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[229]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[229]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[230]~FF  (.D(\test_module/n33 [230]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[230])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[230]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[230]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[230]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[230]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[230]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[230]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[230]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[231]~FF  (.D(\test_module/n33 [231]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[231])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[231]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[231]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[231]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[231]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[231]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[231]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[231]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[232]~FF  (.D(\test_module/n33 [232]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[232])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[232]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[232]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[232]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[232]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[232]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[232]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[232]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[233]~FF  (.D(\test_module/n33 [233]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[233])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[233]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[233]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[233]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[233]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[233]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[233]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[233]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[234]~FF  (.D(\test_module/n33 [234]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[234])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[234]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[234]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[234]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[234]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[234]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[234]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[234]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[235]~FF  (.D(\test_module/n33 [235]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[235])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[235]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[235]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[235]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[235]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[235]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[235]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[235]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[236]~FF  (.D(\test_module/n33 [236]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[236])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[236]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[236]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[236]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[236]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[236]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[236]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[236]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[237]~FF  (.D(\test_module/n33 [237]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[237])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[237]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[237]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[237]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[237]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[237]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[237]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[237]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[238]~FF  (.D(\test_module/n33 [238]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[238])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[238]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[238]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[238]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[238]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[238]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[238]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[238]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[239]~FF  (.D(\test_module/n33 [239]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[239])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[239]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[239]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[239]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[239]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[239]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[239]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[239]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[240]~FF  (.D(\test_module/n33 [240]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[240])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[240]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[240]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[240]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[240]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[240]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[240]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[240]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[241]~FF  (.D(\test_module/n33 [241]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[241])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[241]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[241]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[241]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[241]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[241]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[241]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[241]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[242]~FF  (.D(\test_module/n33 [242]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[242])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[242]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[242]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[242]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[242]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[242]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[242]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[242]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[243]~FF  (.D(\test_module/n33 [243]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[243])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[243]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[243]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[243]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[243]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[243]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[243]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[243]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[244]~FF  (.D(\test_module/n33 [244]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[244])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[244]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[244]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[244]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[244]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[244]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[244]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[244]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[245]~FF  (.D(\test_module/n33 [245]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[245])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[245]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[245]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[245]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[245]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[245]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[245]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[245]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[246]~FF  (.D(\test_module/n33 [246]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[246])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[246]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[246]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[246]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[246]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[246]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[246]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[246]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[247]~FF  (.D(\test_module/n33 [247]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[247])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[247]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[247]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[247]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[247]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[247]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[247]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[247]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[248]~FF  (.D(\test_module/n33 [248]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[248])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[248]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[248]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[248]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[248]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[248]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[248]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[248]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[249]~FF  (.D(\test_module/n33 [249]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[249])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[249]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[249]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[249]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[249]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[249]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[249]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[249]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[250]~FF  (.D(\test_module/n33 [250]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[250])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[250]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[250]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[250]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[250]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[250]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[250]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[250]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[251]~FF  (.D(\test_module/n33 [251]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[251])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[251]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[251]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[251]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[251]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[251]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[251]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[251]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[252]~FF  (.D(\test_module/n33 [252]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[252])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[252]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[252]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[252]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[252]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[252]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[252]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[252]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[253]~FF  (.D(\test_module/n33 [253]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[253])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[253]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[253]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[253]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[253]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[253]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[253]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[253]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[254]~FF  (.D(\test_module/n33 [254]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[254])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[254]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[254]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[254]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[254]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[254]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[254]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[254]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_pllBr0_reg[255]~FF  (.D(\test_module/n33 [255]), .CE(\~test_module/equal_8/n41 ), 
           .CLK(\clk_0~O ), .SR(i_reg_rstn), .Q(o_pllBr0_reg[255])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(24)
    defparam \o_pllBr0_reg[255]~FF .CLK_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[255]~FF .CE_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[255]~FF .SR_POLARITY = 1'b0;
    defparam \o_pllBr0_reg[255]~FF .D_POLARITY = 1'b1;
    defparam \o_pllBr0_reg[255]~FF .SR_SYNC = 1'b0;
    defparam \o_pllBr0_reg[255]~FF .SR_VALUE = 1'b0;
    defparam \o_pllBr0_reg[255]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/internal_reg_r0[0]~FF  (.D(\debug_inst/edb_user_dr [70]), 
           .CE(\debug_inst/vio0/vio_core_inst/n251 ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1395)
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[0]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[0]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[0]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[0]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[0]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[0]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/bit_count[0]~FF  (.D(\debug_inst/vio0/vio_core_inst/n422 [0]), 
           .CE(ceg_net8), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/bit_count [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1429)
    defparam \debug_inst/vio0/vio_core_inst/bit_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[0]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[0]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[0]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[0]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/word_count[0]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_word_counter [0]), 
           .CE(\debug_inst/vio0/vio_core_inst/word_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/word_count [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1447)
    defparam \debug_inst/vio0/vio_core_inst/word_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[0]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[0]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[0]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[0]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_out_shift_reg[0]~FF  (.D(\debug_inst/vio0/vio_core_inst/n546 [0]), 
           .CE(ceg_net11), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[0]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/module_state[0]~FF  (.D(\debug_inst/vio0/vio_core_inst/module_next_state [0]), 
           .CE(1'b1), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/module_state [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1502)
    defparam \debug_inst/vio0/vio_core_inst/module_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/module_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/module_state[0]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/module_state[0]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/module_state[0]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/module_state[0]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/module_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_from_biu[1]~FF  (.D(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [1]), 
           .CE(\debug_inst/vio0/vio_core_inst/n2907 ), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/data_from_biu [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1842)
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[1]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[1]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[1]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[1]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[1]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_from_biu[0]~FF  (.D(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [0]), 
           .CE(\debug_inst/vio0/vio_core_inst/n2907 ), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/data_from_biu [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1842)
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[0]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[0]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[0]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[0]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[0]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/internal_reg_r0[1]~FF  (.D(\debug_inst/edb_user_dr [71]), 
           .CE(\debug_inst/vio0/vio_core_inst/n251 ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1395)
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[1]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[1]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[1]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[1]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[1]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[1]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_from_biu[15]~FF  (.D(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [15]), 
           .CE(\debug_inst/vio0/vio_core_inst/n2907 ), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/data_from_biu [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1842)
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[15]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[15]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[15]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[15]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[15]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[15]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_from_biu[14]~FF  (.D(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [14]), 
           .CE(\debug_inst/vio0/vio_core_inst/n2907 ), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/data_from_biu [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1842)
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[14]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[14]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[14]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[14]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[14]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[14]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_from_biu[13]~FF  (.D(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [13]), 
           .CE(\debug_inst/vio0/vio_core_inst/n2907 ), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/data_from_biu [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1842)
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[13]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[13]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[13]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[13]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[13]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[13]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_from_biu[12]~FF  (.D(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [12]), 
           .CE(\debug_inst/vio0/vio_core_inst/n2907 ), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/data_from_biu [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1842)
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[12]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[12]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[12]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[12]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[12]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[12]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_from_biu[11]~FF  (.D(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [11]), 
           .CE(\debug_inst/vio0/vio_core_inst/n2907 ), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/data_from_biu [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1842)
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[11]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[11]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[11]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[11]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[11]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[11]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_from_biu[10]~FF  (.D(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [10]), 
           .CE(\debug_inst/vio0/vio_core_inst/n2907 ), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/data_from_biu [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1842)
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[10]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[10]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[10]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[10]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[10]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[10]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_from_biu[9]~FF  (.D(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [9]), 
           .CE(\debug_inst/vio0/vio_core_inst/n2907 ), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/data_from_biu [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1842)
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[9]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[9]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[9]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[9]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[9]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_from_biu[8]~FF  (.D(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [8]), 
           .CE(\debug_inst/vio0/vio_core_inst/n2907 ), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/data_from_biu [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1842)
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[8]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[8]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[8]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[8]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[8]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_from_biu[7]~FF  (.D(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [7]), 
           .CE(\debug_inst/vio0/vio_core_inst/n2907 ), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/data_from_biu [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1842)
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[7]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[7]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[7]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[7]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[7]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_from_biu[6]~FF  (.D(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [6]), 
           .CE(\debug_inst/vio0/vio_core_inst/n2907 ), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/data_from_biu [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1842)
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[6]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[6]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[6]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[6]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[6]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_from_biu[5]~FF  (.D(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [5]), 
           .CE(\debug_inst/vio0/vio_core_inst/n2907 ), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/data_from_biu [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1842)
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[5]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[5]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[5]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[5]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[5]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_from_biu[4]~FF  (.D(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [4]), 
           .CE(\debug_inst/vio0/vio_core_inst/n2907 ), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/data_from_biu [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1842)
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[4]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[4]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[4]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[4]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[4]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_from_biu[3]~FF  (.D(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [3]), 
           .CE(\debug_inst/vio0/vio_core_inst/n2907 ), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/data_from_biu [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1842)
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[3]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[3]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[3]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[3]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[3]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_from_biu[2]~FF  (.D(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [2]), 
           .CE(\debug_inst/vio0/vio_core_inst/n2907 ), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/data_from_biu [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1842)
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[2]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[2]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[2]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[2]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[2]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_from_biu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[31]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [31]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[31]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[31]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[31]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[31]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[31]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[31]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[30]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [30]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[30]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[30]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[30]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[30]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[30]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[30]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[29]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [29]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[29]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[29]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[29]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[29]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[29]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[29]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[28]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [28]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[28]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[28]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[28]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[28]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[28]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[28]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[27]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [27]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[27]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[27]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[27]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[27]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[27]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[27]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[26]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [26]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[26]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[26]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[26]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[26]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[26]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[26]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[25]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [25]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[25]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[25]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[25]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[25]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[25]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[25]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[24]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [24]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[24]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[24]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[24]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[24]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[24]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[24]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[23]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [23]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[23]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[23]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[23]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[23]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[23]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[23]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[22]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [22]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[22]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[22]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[22]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[22]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[22]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[22]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[21]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [21]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[21]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[21]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[21]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[21]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[21]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[21]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[20]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [20]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[20]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[20]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[20]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[20]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[20]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[20]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[19]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [19]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[19]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[19]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[19]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[19]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[19]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[19]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[18]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [18]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[18]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[18]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[18]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[18]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[18]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[18]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[17]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [17]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[17]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[17]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[17]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[17]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[17]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[17]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[16]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [16]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[16]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[16]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[16]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[16]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[16]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[16]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[15]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [15]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[15]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[15]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[15]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[15]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[15]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[15]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[14]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [14]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[14]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[14]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[14]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[14]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[14]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[14]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[13]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [13]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[13]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[13]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[13]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[13]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[13]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[13]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[12]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [12]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[12]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[12]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[12]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[12]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[12]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[12]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[11]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [11]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[11]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[11]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[11]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[11]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[11]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[11]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[10]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [10]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[10]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[10]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[10]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[10]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[10]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[10]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[9]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [9]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[9]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[9]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[9]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[9]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[9]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[9]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[8]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [8]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[8]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[8]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[8]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[8]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[8]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[8]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[7]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [7]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[7]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[7]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[7]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[7]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[7]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[7]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[6]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [6]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[6]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[6]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[6]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[6]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[6]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[6]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[5]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [5]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[5]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[5]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[5]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[5]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[5]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[5]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[4]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [4]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[4]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[4]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[4]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[4]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[4]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[4]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[3]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [3]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[3]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[3]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[3]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[3]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[3]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[3]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[2]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [2]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[2]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[2]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[2]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[2]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[2]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[2]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[1]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [1]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[1]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[1]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[1]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[1]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[1]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[1]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/crc_data_out[0]~FF  (.D(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [0]), 
           .CE(ceg_net16), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/crc_data_out [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[0]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[0]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[0]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[0]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[0]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[0]~FF .SR_VALUE = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/crc_data_out[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/module_state[3]~FF  (.D(\debug_inst/vio0/vio_core_inst/module_next_state [3]), 
           .CE(1'b1), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/module_state [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1502)
    defparam \debug_inst/vio0/vio_core_inst/module_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/module_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/module_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/module_state[3]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/module_state[3]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/module_state[3]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/module_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/module_state[2]~FF  (.D(\debug_inst/vio0/vio_core_inst/module_next_state [2]), 
           .CE(1'b1), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/module_state [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1502)
    defparam \debug_inst/vio0/vio_core_inst/module_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/module_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/module_state[2]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/module_state[2]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/module_state[2]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/module_state[2]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/module_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/module_state[1]~FF  (.D(\debug_inst/vio0/vio_core_inst/module_next_state [1]), 
           .CE(1'b1), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/module_state [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1502)
    defparam \debug_inst/vio0/vio_core_inst/module_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/module_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/module_state[1]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/module_state[1]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/module_state[1]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/module_state[1]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/module_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_out_shift_reg[15]~FF  (.D(\debug_inst/vio0/vio_core_inst/n546 [15]), 
           .CE(ceg_net11), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[15]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_out_shift_reg[14]~FF  (.D(\debug_inst/vio0/vio_core_inst/n546 [14]), 
           .CE(ceg_net11), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[14]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[14]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[14]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[14]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[14]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[14]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_out_shift_reg[13]~FF  (.D(\debug_inst/vio0/vio_core_inst/n546 [13]), 
           .CE(ceg_net11), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[13]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[13]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[13]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[13]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[13]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[13]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_out_shift_reg[12]~FF  (.D(\debug_inst/vio0/vio_core_inst/n546 [12]), 
           .CE(ceg_net11), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[12]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[12]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[12]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[12]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[12]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[12]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_out_shift_reg[11]~FF  (.D(\debug_inst/vio0/vio_core_inst/n546 [11]), 
           .CE(ceg_net11), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[11]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[11]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[11]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[11]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[11]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[11]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_out_shift_reg[10]~FF  (.D(\debug_inst/vio0/vio_core_inst/n546 [10]), 
           .CE(ceg_net11), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[10]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[10]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[10]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[10]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[10]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[10]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_out_shift_reg[9]~FF  (.D(\debug_inst/vio0/vio_core_inst/n546 [9]), 
           .CE(ceg_net11), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[9]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[9]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[9]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[9]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[9]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[9]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_out_shift_reg[8]~FF  (.D(\debug_inst/vio0/vio_core_inst/n546 [8]), 
           .CE(ceg_net11), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[8]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[8]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[8]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[8]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[8]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[8]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_out_shift_reg[7]~FF  (.D(\debug_inst/vio0/vio_core_inst/n546 [7]), 
           .CE(ceg_net11), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[7]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[7]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[7]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_out_shift_reg[6]~FF  (.D(\debug_inst/vio0/vio_core_inst/n546 [6]), 
           .CE(ceg_net11), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[6]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[6]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[6]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_out_shift_reg[5]~FF  (.D(\debug_inst/vio0/vio_core_inst/n546 [5]), 
           .CE(ceg_net11), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[5]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[5]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[5]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_out_shift_reg[4]~FF  (.D(\debug_inst/vio0/vio_core_inst/n546 [4]), 
           .CE(ceg_net11), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[4]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[4]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_out_shift_reg[3]~FF  (.D(\debug_inst/vio0/vio_core_inst/n546 [3]), 
           .CE(ceg_net11), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[3]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_out_shift_reg[2]~FF  (.D(\debug_inst/vio0/vio_core_inst/n546 [2]), 
           .CE(ceg_net11), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[2]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/data_out_shift_reg[1]~FF  (.D(\debug_inst/vio0/vio_core_inst/n546 [1]), 
           .CE(ceg_net11), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[1]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/data_out_shift_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/word_count[15]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_word_counter [15]), 
           .CE(\debug_inst/vio0/vio_core_inst/word_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/word_count [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1447)
    defparam \debug_inst/vio0/vio_core_inst/word_count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[15]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[15]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[15]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[15]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[15]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/word_count[14]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_word_counter [14]), 
           .CE(\debug_inst/vio0/vio_core_inst/word_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/word_count [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1447)
    defparam \debug_inst/vio0/vio_core_inst/word_count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[14]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[14]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[14]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[14]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[14]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/word_count[13]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_word_counter [13]), 
           .CE(\debug_inst/vio0/vio_core_inst/word_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/word_count [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1447)
    defparam \debug_inst/vio0/vio_core_inst/word_count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[13]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[13]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[13]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[13]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[13]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/word_count[12]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_word_counter [12]), 
           .CE(\debug_inst/vio0/vio_core_inst/word_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/word_count [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1447)
    defparam \debug_inst/vio0/vio_core_inst/word_count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[12]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[12]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[12]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[12]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[12]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/word_count[11]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_word_counter [11]), 
           .CE(\debug_inst/vio0/vio_core_inst/word_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/word_count [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1447)
    defparam \debug_inst/vio0/vio_core_inst/word_count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[11]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[11]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[11]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[11]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[11]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/word_count[10]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_word_counter [10]), 
           .CE(\debug_inst/vio0/vio_core_inst/word_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/word_count [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1447)
    defparam \debug_inst/vio0/vio_core_inst/word_count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[10]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[10]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[10]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[10]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[10]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/word_count[9]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_word_counter [9]), 
           .CE(\debug_inst/vio0/vio_core_inst/word_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/word_count [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1447)
    defparam \debug_inst/vio0/vio_core_inst/word_count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[9]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[9]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[9]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[9]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[9]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/word_count[8]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_word_counter [8]), 
           .CE(\debug_inst/vio0/vio_core_inst/word_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/word_count [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1447)
    defparam \debug_inst/vio0/vio_core_inst/word_count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[8]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[8]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[8]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[8]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[8]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/word_count[7]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_word_counter [7]), 
           .CE(\debug_inst/vio0/vio_core_inst/word_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/word_count [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1447)
    defparam \debug_inst/vio0/vio_core_inst/word_count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[7]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[7]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[7]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[7]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[7]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/word_count[6]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_word_counter [6]), 
           .CE(\debug_inst/vio0/vio_core_inst/word_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/word_count [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1447)
    defparam \debug_inst/vio0/vio_core_inst/word_count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[6]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[6]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[6]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[6]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[6]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/word_count[5]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_word_counter [5]), 
           .CE(\debug_inst/vio0/vio_core_inst/word_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/word_count [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1447)
    defparam \debug_inst/vio0/vio_core_inst/word_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[5]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[5]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[5]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[5]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/word_count[4]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_word_counter [4]), 
           .CE(\debug_inst/vio0/vio_core_inst/word_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/word_count [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1447)
    defparam \debug_inst/vio0/vio_core_inst/word_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[4]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[4]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[4]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[4]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/word_count[3]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_word_counter [3]), 
           .CE(\debug_inst/vio0/vio_core_inst/word_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/word_count [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1447)
    defparam \debug_inst/vio0/vio_core_inst/word_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[3]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[3]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[3]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[3]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/word_count[2]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_word_counter [2]), 
           .CE(\debug_inst/vio0/vio_core_inst/word_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/word_count [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1447)
    defparam \debug_inst/vio0/vio_core_inst/word_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[2]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[2]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[2]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[2]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/word_count[1]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_word_counter [1]), 
           .CE(\debug_inst/vio0/vio_core_inst/word_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/word_count [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1447)
    defparam \debug_inst/vio0/vio_core_inst/word_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[1]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[1]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/word_count[1]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[1]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/word_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/bit_count[5]~FF  (.D(\debug_inst/vio0/vio_core_inst/n422 [5]), 
           .CE(ceg_net8), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/bit_count [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1429)
    defparam \debug_inst/vio0/vio_core_inst/bit_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[5]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[5]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[5]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[5]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/bit_count[4]~FF  (.D(\debug_inst/vio0/vio_core_inst/n422 [4]), 
           .CE(ceg_net8), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/bit_count [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1429)
    defparam \debug_inst/vio0/vio_core_inst/bit_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[4]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[4]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[4]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[4]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/bit_count[3]~FF  (.D(\debug_inst/vio0/vio_core_inst/n422 [3]), 
           .CE(ceg_net8), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/bit_count [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1429)
    defparam \debug_inst/vio0/vio_core_inst/bit_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[3]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[3]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[3]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[3]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/bit_count[2]~FF  (.D(\debug_inst/vio0/vio_core_inst/n422 [2]), 
           .CE(ceg_net8), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/bit_count [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1429)
    defparam \debug_inst/vio0/vio_core_inst/bit_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[2]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[2]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[2]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[2]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/bit_count[1]~FF  (.D(\debug_inst/vio0/vio_core_inst/n422 [1]), 
           .CE(ceg_net8), .CLK(\bscan_TCK~O ), .SR(\debug_inst/edb_soft_reset ), 
           .Q(\debug_inst/vio0/vio_core_inst/bit_count [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1429)
    defparam \debug_inst/vio0/vio_core_inst/bit_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[1]~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[1]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[1]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[1]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/bit_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/opcode[2]~FF  (.D(\debug_inst/edb_user_dr [79]), 
           .CE(\debug_inst/vio0/vio_core_inst/op_reg_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/opcode [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1420)
    defparam \debug_inst/vio0/vio_core_inst/opcode[2]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/opcode[2]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/opcode[2]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/opcode[2]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/opcode[2]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/opcode[2]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/opcode[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/opcode[1]~FF  (.D(\debug_inst/edb_user_dr [78]), 
           .CE(\debug_inst/vio0/vio_core_inst/op_reg_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/opcode [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1420)
    defparam \debug_inst/vio0/vio_core_inst/opcode[1]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/opcode[1]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/opcode[1]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/opcode[1]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/opcode[1]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/opcode[1]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/opcode[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/address_counter[5]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_addr_counter [5]), 
           .CE(\debug_inst/vio0/vio_core_inst/addr_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/address_counter [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1410)
    defparam \debug_inst/vio0/vio_core_inst/address_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[5]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[5]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/address_counter[4]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_addr_counter [4]), 
           .CE(\debug_inst/vio0/vio_core_inst/addr_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/address_counter [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1410)
    defparam \debug_inst/vio0/vio_core_inst/address_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[4]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[4]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/address_counter[3]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_addr_counter [3]), 
           .CE(\debug_inst/vio0/vio_core_inst/addr_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/address_counter [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1410)
    defparam \debug_inst/vio0/vio_core_inst/address_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[3]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[3]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/address_counter[2]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_addr_counter [2]), 
           .CE(\debug_inst/vio0/vio_core_inst/addr_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/address_counter [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1410)
    defparam \debug_inst/vio0/vio_core_inst/address_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[2]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[2]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/address_counter[1]~FF  (.D(\debug_inst/vio0/vio_core_inst/data_to_addr_counter [1]), 
           .CE(\debug_inst/vio0/vio_core_inst/addr_ct_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/address_counter [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1410)
    defparam \debug_inst/vio0/vio_core_inst/address_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[1]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[1]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[1]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/address_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/internal_reg_r0[2]~FF  (.D(\debug_inst/edb_user_dr [72]), 
           .CE(\debug_inst/vio0/vio_core_inst/n251 ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1395)
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[2]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[2]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[2]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[2]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[2]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[2]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/internal_reg_r0[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/commit_sync1~FF  (.D(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [0]), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/commit_sync1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1849)
    defparam \debug_inst/vio0/vio_core_inst/commit_sync1~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/commit_sync1~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/commit_sync1~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/commit_sync1~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/commit_sync1~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/commit_sync1~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/commit_sync1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/commit_sync2~FF  (.D(\debug_inst/vio0/vio_core_inst/commit_sync1 ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/commit_sync2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1849)
    defparam \debug_inst/vio0/vio_core_inst/commit_sync2~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/commit_sync2~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/commit_sync2~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/commit_sync2~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/commit_sync2~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/commit_sync2~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/commit_sync2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i_reg_rstn~FF  (.D(\debug_inst/vio0/vio_core_inst/probe_out_sync [0]), 
           .CE(\debug_inst/vio0/vio_core_inst/commit_sync2 ), .CLK(\clk_0~O ), 
           .SR(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [1]), .Q(i_reg_rstn)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1857)
    defparam \i_reg_rstn~FF .CLK_POLARITY = 1'b1;
    defparam \i_reg_rstn~FF .CE_POLARITY = 1'b1;
    defparam \i_reg_rstn~FF .SR_POLARITY = 1'b1;
    defparam \i_reg_rstn~FF .D_POLARITY = 1'b1;
    defparam \i_reg_rstn~FF .SR_SYNC = 1'b0;
    defparam \i_reg_rstn~FF .SR_VALUE = 1'b0;
    defparam \i_reg_rstn~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_out_sync[0]~FF  (.D(\debug_inst/edb_user_dr [67]), 
           .CE(\debug_inst/vio0/vio_core_inst/n2952 ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [1]), .Q(\debug_inst/vio0/vio_core_inst/probe_out_sync [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1868)
    defparam \debug_inst/vio0/vio_core_inst/probe_out_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_out_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_out_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_out_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_out_sync[0]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_out_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_out_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/internal_register_select[0]~FF  (.D(\debug_inst/edb_user_dr [73]), 
           .CE(\debug_inst/vio0/vio_core_inst/regsel_ld_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/internal_register_select [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1351)
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[0]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[0]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[0]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[0]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[0]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[0]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[0]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[0]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[0]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[0].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[1]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[1]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[1]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[1]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[1].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[2]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[2]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[2]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[2]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[2]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[2]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[2]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[2]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[2].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[3]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[3]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[3]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[3]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[3]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[3]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[3]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[3]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[3].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[4]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[4]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[4].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[5]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[5]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[5].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[6]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[6]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[6].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[7]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[7]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[7].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[8]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[8]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[8].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[9]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[9]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[9]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[9]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[9]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[9]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[9]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[9]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[9].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[10]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[10]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[10]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[10]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[10]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[10]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[10]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[10]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[10].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[11]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[11]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[11]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[11]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[11]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[11]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[11]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[11]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[11].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[12]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[12]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[12]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[12]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[12]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[12]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[12]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[12]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[12].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[13]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[13]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[13]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[13]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[13]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[13]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[13]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[13]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[13].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[14]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[14]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[14]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[14]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[14]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[14]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[14]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[14]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[14].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[15]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[15]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[15]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[15]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[15]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[15]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[15]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[15]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[15].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[16]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[16]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[16]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[16]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[16]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[16]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[16]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[16]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[16].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[17]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[17]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[17]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[17]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[17]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[17]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[17]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[17]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[17].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[18]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[18]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[18]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[18]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[18]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[18]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[18]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[18]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[18].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[19]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[19]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[19]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[19]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[19]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[19]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[19]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[19]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[19].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[20]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[20]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[20]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[20]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[20]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[20]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[20]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[20]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[20].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[21]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[21]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[21]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[21]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[21]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[21]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[21]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[21]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[21].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[22]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[22]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[22]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[22]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[22]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[22]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[22]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[22]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[22].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[23]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[23]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[23]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[23]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[23]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[23]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[23]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[23]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[23].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[24]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[24]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[24]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[24]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[24]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[24]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[24]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[24]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[24].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[25]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[25]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[25]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[25]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[25]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[25]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[25]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[25]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[25].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[26]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[26]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[26]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[26]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[26]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[26]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[26]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[26]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[26].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[27]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[27]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[27]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[27]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[27]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[27]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[27]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[27]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[27].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[28]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[28]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[28]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[28]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[28]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[28]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[28]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[28]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[28].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[29]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[29]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[29]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[29]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[29]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[29]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[29]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[29]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[29].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[30]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[30]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[30]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[30]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[30]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[30]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[30]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[30]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[30].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[31]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[31]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[31]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[31]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[31]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[31]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[31]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[31]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[31].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[32]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[32]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[32]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[32]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[32]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[32]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[32]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[32]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[32].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[33]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[33]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[33]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[33]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[33]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[33]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[33]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[33]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[33].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[34]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[34]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[34]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[34]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[34]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[34]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[34]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[34]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[34].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[35]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[35]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[35]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[35]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[35]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[35]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[35]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[35]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[35].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[36]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[36]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[36]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[36]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[36]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[36]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[36]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[36]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[36].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[37]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[37]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[37]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[37]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[37]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[37]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[37]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[37]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[37].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[38]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[38]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[38]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[38]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[38]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[38]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[38]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[38]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[38].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[39]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[39]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[39]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[39]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[39]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[39]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[39]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[39]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[39].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[40]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[40]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[40]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[40]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[40]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[40]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[40]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[40]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[40].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[41]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[41]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[41]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[41]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[41]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[41]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[41]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[41]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[41].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[42]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[42]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[42]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[42]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[42]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[42]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[42]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[42]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[42].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[43]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[43]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[43]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[43]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[43]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[43]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[43]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[43]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[43].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[44]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[44]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[44]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[44]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[44]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[44]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[44]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[44]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[44].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[45]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[45]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[45]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[45]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[45]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[45]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[45]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[45]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[45].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[46]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[46]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[46]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[46]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[46]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[46]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[46]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[46]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[46].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[47]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[47]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[47]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[47]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[47]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[47]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[47]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[47]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[47].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[48]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[48]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[48]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[48]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[48]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[48]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[48]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[48]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[48].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[49]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[49]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[49]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[49]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[49]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[49]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[49]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[49]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[49].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[50]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[50]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[50]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[50]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[50]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[50]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[50]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[50]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[50].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[51]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[51]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[51]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[51]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[51]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[51]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[51]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[51]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[51].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[52]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[52]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[52]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[52]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[52]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[52]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[52]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[52]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[52].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[53]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[53]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[53]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[53]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[53]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[53]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[53]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[53]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[53].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[54]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[54]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[54]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[54]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[54]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[54]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[54]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[54]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[54].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[55]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[55]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[55]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[55]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[55]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[55]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[55]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[55]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[55].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[56]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[56]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[56]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[56]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[56]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[56]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[56]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[56]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[56].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[57]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[57]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[57]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[57]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[57]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[57]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[57]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[57]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[57].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[58]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[58]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[58]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[58]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[58]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[58]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[58]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[58]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[58].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[59]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[59]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[59]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[59]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[59]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[59]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[59]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[59]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[59].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[60]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [60])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[60]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[60]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[60]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[60]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[60]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[60]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[60]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[60].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[61]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [61])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[61]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[61]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[61]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[61]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[61]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[61]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[61]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[61].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[62]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [62])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[62]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[62]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[62]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[62]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[62]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[62]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[62]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[62].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[63]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[63]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[63]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[63]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[63]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[63]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[63]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[63]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[63].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[64]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [64])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[64]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[64]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[64]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[64]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[64]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[64]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[64]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[64].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[65]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [65])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[65]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[65]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[65]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[65]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[65]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[65]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[65]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[65].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[66]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [66])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[66]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[66]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[66]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[66]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[66]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[66]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[66]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[66].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[67]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [67])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[67]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[67]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[67]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[67]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[67]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[67]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[67]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[67].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[68]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [68])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[68]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[68]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[68]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[68]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[68]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[68]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[68]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[68].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[69]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [69])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[69]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[69]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[69]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[69]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[69]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[69]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[69]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[69].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[70]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [70])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[70]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[70]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[70]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[70]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[70]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[70]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[70]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[70].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[71]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [71])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[71]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[71]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[71]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[71]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[71]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[71]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[71]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[71].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[72]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [72])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[72]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[72]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[72]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[72]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[72]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[72]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[72]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[72].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[73]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [73])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[73]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[73]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[73]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[73]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[73]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[73]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[73]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[73].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[74]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [74])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[74]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[74]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[74]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[74]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[74]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[74]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[74]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[74].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[75]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [75])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[75]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[75]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[75]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[75]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[75]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[75]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[75]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[75].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[76]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [76])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[76]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[76]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[76]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[76]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[76]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[76]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[76]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[76].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[77]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [77])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[77]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[77]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[77]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[77]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[77]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[77]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[77]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[77].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[78]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [78])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[78]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[78]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[78]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[78]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[78]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[78]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[78]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[78].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[79]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [79])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[79]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[79]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[79]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[79]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[79]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[79]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[79]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[79].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[80]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [80])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[80]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[80]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[80]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[80]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[80]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[80]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[80]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[80].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[81]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [81])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[81]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[81]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[81]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[81]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[81]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[81]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[81]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[81].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[82]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [82])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[82]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[82]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[82]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[82]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[82]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[82]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[82]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[82].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[83]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [83])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[83]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[83]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[83]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[83]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[83]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[83]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[83]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[83].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[84]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [84])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[84]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[84]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[84]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[84]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[84]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[84]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[84]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[84].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[85]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [85])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[85]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[85]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[85]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[85]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[85]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[85]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[85]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[85].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[86]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [86])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[86]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[86]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[86]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[86]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[86]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[86]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[86]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[86].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[87]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [87])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[87]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[87]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[87]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[87]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[87]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[87]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[87]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[87].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[88]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [88])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[88]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[88]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[88]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[88]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[88]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[88]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[88]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[88].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[89]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [89])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[89]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[89]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[89]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[89]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[89]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[89]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[89]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[89].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[90]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [90])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[90]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[90]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[90]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[90]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[90]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[90]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[90]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[90].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[91]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [91])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[91]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[91]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[91]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[91]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[91]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[91]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[91]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[91].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[92]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [92])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[92]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[92]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[92]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[92]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[92]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[92]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[92]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[92].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[93]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [93])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[93]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[93]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[93]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[93]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[93]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[93]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[93]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[93].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[94]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [94])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[94]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[94]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[94]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[94]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[94]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[94]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[94]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[94].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[95]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [95])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[95]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[95]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[95]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[95]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[95]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[95]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[95]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[95].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[96]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [96])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[96]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[96]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[96]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[96]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[96]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[96]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[96]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[96].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[97]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [97])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[97]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[97]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[97]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[97]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[97]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[97]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[97]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[97].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[98]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [98])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[98]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[98]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[98]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[98]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[98]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[98]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[98]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[98].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[99]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [99])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[99]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[99]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[99]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[99]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[99]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[99]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[99]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[99].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[100]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [100])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[100]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[100]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[100]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[100]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[100]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[100]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[100]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[100].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[101]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [101])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[101]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[101]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[101]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[101]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[101]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[101]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[101]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[101].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[102]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [102])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[102]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[102]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[102]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[102]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[102]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[102]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[102]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[102].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[103]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [103])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[103]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[103]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[103]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[103]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[103]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[103]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[103]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[103].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[104]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [104])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[104]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[104]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[104]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[104]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[104]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[104]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[104]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[104].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[105]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [105])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[105]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[105]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[105]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[105]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[105]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[105]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[105]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[105].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[106]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [106])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[106]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[106]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[106]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[106]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[106]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[106]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[106]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[106].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[107]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [107])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[107]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[107]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[107]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[107]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[107]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[107]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[107]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[107].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[108]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [108])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[108]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[108]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[108]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[108]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[108]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[108]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[108]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[108].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[109]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [109])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[109]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[109]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[109]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[109]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[109]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[109]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[109]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[109].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[110]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [110])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[110]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[110]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[110]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[110]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[110]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[110]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[110]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[110].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[111]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [111])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[111]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[111]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[111]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[111]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[111]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[111]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[111]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[111].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[112]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [112])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[112]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[112]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[112]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[112]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[112]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[112]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[112]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[112].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[113]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [113])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[113]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[113]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[113]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[113]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[113]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[113]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[113]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[113].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[114]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [114])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[114]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[114]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[114]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[114]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[114]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[114]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[114]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[114].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[115]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [115])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[115]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[115]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[115]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[115]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[115]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[115]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[115]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[115].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[116]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [116])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[116]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[116]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[116]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[116]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[116]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[116]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[116]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[116].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[117]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [117])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[117]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[117]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[117]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[117]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[117]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[117]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[117]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[117].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[118]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [118])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[118]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[118]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[118]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[118]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[118]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[118]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[118]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[118].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[119]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [119])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[119]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[119]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[119]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[119]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[119]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[119]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[119]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[119].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[120]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [120])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[120]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[120]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[120]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[120]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[120]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[120]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[120]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[120]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[120].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[121]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [121])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[121]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[121]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[121]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[121]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[121]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[121]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[121]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[121]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[121].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[122]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [122])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[122]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[122]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[122]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[122]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[122]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[122]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[122]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[122]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[122].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[123]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [123])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[123]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[123]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[123]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[123]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[123]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[123]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[123]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[123]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[123].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[124]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [124])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[124]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[124]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[124]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[124]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[124]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[124]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[124]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[124]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[124].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[125]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [125])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[125]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[125]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[125]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[125]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[125]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[125]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[125]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[125]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[125].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[126]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [126])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[126]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[126]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[126]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[126]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[126]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[126]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[126]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[126]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[126].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[127]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [127])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[127]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[127]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[127]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[127]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[127]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[127]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[127]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[127]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[127].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[128]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [128])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[128]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[128]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[128]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[128]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[128]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[128]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[128]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[128]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[128].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[129]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [129])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[129]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[129]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[129]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[129]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[129]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[129]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[129]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[129]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[129].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[130]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [130])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[130]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[130]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[130]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[130]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[130]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[130]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[130]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[130]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[130].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[131]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [131])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[131]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[131]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[131]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[131]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[131]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[131]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[131]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[131]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[131].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[132]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [132])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[132]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[132]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[132]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[132]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[132]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[132]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[132]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[132]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[132].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[133]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [133])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[133]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[133]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[133]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[133]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[133]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[133]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[133]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[133]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[133].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[134]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [134])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[134]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[134]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[134]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[134]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[134]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[134]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[134]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[134]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[134].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[135]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [135])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[135]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[135]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[135]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[135]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[135]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[135]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[135]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[135]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[135].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[136]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [136])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[136]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[136]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[136]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[136]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[136]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[136]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[136]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[136]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[136].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[137]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [137])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[137]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[137]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[137]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[137]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[137]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[137]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[137]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[137]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[137].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[138]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [138])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[138]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[138]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[138]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[138]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[138]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[138]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[138]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[138]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[138].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[139]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [139])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[139]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[139]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[139]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[139]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[139]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[139]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[139]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[139]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[139].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[140]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [140])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[140]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[140]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[140]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[140]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[140]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[140]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[140]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[140]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[140].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[141]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [141])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[141]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[141]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[141]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[141]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[141]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[141]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[141]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[141]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[141].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[142]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [142])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[142]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[142]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[142]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[142]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[142]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[142]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[142]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[142]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[142].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[143]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [143])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[143]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[143]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[143]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[143]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[143]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[143]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[143]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[143]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[143].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[144]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [144])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[144]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[144]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[144]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[144]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[144]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[144]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[144]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[144]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[144].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[145]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [145])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[145]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[145]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[145]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[145]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[145]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[145]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[145]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[145]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[145].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[146]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [146])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[146]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[146]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[146]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[146]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[146]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[146]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[146]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[146]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[146].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[147]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [147])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[147]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[147]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[147]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[147]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[147]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[147]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[147]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[147]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[147].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[148]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [148])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[148]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[148]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[148]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[148]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[148]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[148]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[148]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[148]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[148].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[149]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [149])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[149]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[149]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[149]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[149]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[149]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[149]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[149]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[149]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[149].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[150]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [150])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[150]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[150]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[150]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[150]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[150]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[150]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[150]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[150]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[150].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[151]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [151])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[151]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[151]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[151]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[151]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[151]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[151]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[151]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[151]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[151].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[152]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [152])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[152]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[152]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[152]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[152]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[152]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[152]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[152]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[152]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[152].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[153]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [153])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[153]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[153]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[153]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[153]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[153]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[153]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[153]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[153]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[153].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[154]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [154])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[154]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[154]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[154]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[154]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[154]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[154]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[154]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[154]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[154].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[155]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [155])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[155]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[155]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[155]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[155]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[155]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[155]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[155]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[155]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[155].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[156]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [156])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[156]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[156]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[156]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[156]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[156]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[156]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[156]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[156]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[156].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[157]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [157])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[157]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[157]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[157]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[157]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[157]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[157]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[157]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[157]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[157].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[158]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [158])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[158]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[158]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[158]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[158]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[158]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[158]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[158]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[158]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[158].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[159]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [159])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[159]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[159]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[159]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[159]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[159]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[159]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[159]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[159]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[159].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[160]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [160])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[160]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[160]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[160]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[160]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[160]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[160]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[160]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[160]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[160].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[161]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [161])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[161]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[161]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[161]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[161]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[161]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[161]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[161]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[161]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[161].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[162]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [162])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[162]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[162]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[162]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[162]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[162]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[162]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[162]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[162]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[162].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[163]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [163])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[163]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[163]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[163]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[163]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[163]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[163]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[163]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[163]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[163].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[164]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [164])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[164]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[164]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[164]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[164]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[164]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[164]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[164]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[164]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[164].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[165]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [165])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[165]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[165]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[165]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[165]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[165]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[165]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[165]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[165]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[165].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[166]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [166])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[166]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[166]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[166]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[166]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[166]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[166]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[166]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[166]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[166].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[167]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [167])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[167]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[167]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[167]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[167]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[167]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[167]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[167]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[167]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[167].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[168]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [168])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[168]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[168]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[168]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[168]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[168]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[168]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[168]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[168]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[168].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[169]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [169])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[169]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[169]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[169]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[169]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[169]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[169]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[169]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[169]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[169].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[170]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [170])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[170]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[170]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[170]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[170]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[170]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[170]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[170]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[170]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[170].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[171]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [171])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[171]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[171]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[171]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[171]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[171]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[171]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[171]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[171]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[171].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[172]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [172])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[172]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[172]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[172]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[172]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[172]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[172]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[172]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[172]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[172].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[173]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [173])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[173]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[173]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[173]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[173]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[173]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[173]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[173]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[173]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[173].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[174]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [174])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[174]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[174]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[174]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[174]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[174]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[174]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[174]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[174]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[174].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[175]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [175])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[175]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[175]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[175]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[175]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[175]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[175]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[175]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[175]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[175].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[176]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [176])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[176]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[176]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[176]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[176]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[176]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[176]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[176]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[176]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[176].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[177]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [177])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[177]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[177]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[177]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[177]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[177]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[177]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[177]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[177]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[177].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[178]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [178])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[178]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[178]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[178]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[178]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[178]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[178]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[178]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[178]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[178].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[179]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [179])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[179]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[179]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[179]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[179]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[179]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[179]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[179]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[179]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[179].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[180]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [180])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[180]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[180]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[180]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[180]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[180]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[180]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[180]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[180]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[180].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[181]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [181])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[181]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[181]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[181]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[181]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[181]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[181]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[181]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[181]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[181].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[182]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [182])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[182]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[182]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[182]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[182]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[182]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[182]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[182]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[182]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[182].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[183]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [183])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[183]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[183]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[183]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[183]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[183]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[183]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[183]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[183]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[183].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[184]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [184])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[184]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[184]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[184]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[184]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[184]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[184]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[184]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[184]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[184].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[185]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [185])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[185]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[185]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[185]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[185]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[185]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[185]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[185]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[185]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[185].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[186]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [186])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[186]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[186]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[186]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[186]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[186]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[186]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[186]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[186]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[186].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[187]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [187])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[187]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[187]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[187]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[187]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[187]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[187]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[187]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[187]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[187].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[188]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [188])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[188]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[188]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[188]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[188]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[188]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[188]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[188]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[188]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[188].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[189]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [189])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[189]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[189]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[189]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[189]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[189]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[189]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[189]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[189]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[189].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[190]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [190])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[190]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[190]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[190]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[190]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[190]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[190]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[190]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[190]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[190].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[191]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [191])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[191]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[191]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[191]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[191]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[191]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[191]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[191]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[191]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[191].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[192]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [192])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[192]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[192]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[192]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[192]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[192]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[192]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[192]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[192]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[192].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[193]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [193])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[193]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[193]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[193]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[193]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[193]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[193]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[193]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[193]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[193].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[194]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [194])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[194]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[194]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[194]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[194]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[194]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[194]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[194]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[194]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[194].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[195]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [195])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[195]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[195]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[195]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[195]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[195]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[195]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[195]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[195]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[195].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[196]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [196])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[196]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[196]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[196]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[196]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[196]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[196]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[196]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[196]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[196].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[197]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [197])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[197]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[197]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[197]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[197]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[197]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[197]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[197]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[197]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[197].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[198]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [198])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[198]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[198]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[198]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[198]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[198]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[198]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[198]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[198]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[198].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[199]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [199])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[199]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[199]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[199]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[199]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[199]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[199]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[199]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[199]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[199].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[200]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [200])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[200]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[200]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[200]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[200]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[200]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[200]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[200]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[200]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[200].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[201]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [201])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[201]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[201]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[201]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[201]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[201]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[201]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[201]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[201]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[201].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[202]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [202])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[202]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[202]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[202]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[202]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[202]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[202]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[202]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[202]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[202].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[203]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [203])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[203]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[203]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[203]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[203]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[203]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[203]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[203]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[203]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[203].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[204]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [204])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[204]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[204]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[204]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[204]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[204]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[204]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[204]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[204]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[204].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[205]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [205])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[205]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[205]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[205]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[205]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[205]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[205]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[205]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[205]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[205].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[206]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [206])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[206]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[206]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[206]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[206]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[206]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[206]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[206]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[206]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[206].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[207]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [207])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[207]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[207]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[207]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[207]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[207]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[207]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[207]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[207]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[207].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[208]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [208])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[208]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[208]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[208]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[208]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[208]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[208]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[208]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[208]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[208].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[209]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [209])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[209]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[209]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[209]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[209]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[209]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[209]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[209]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[209]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[209].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[210]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [210])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[210]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[210]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[210]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[210]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[210]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[210]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[210]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[210]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[210].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[211]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [211])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[211]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[211]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[211]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[211]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[211]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[211]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[211]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[211]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[211].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[212]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [212])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[212]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[212]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[212]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[212]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[212]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[212]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[212]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[212]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[212].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[213]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [213])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[213]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[213]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[213]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[213]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[213]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[213]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[213]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[213]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[213].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[214]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [214])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[214]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[214]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[214]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[214]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[214]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[214]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[214]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[214]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[214].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[215]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [215])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[215]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[215]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[215]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[215]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[215]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[215]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[215]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[215]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[215].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[216]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [216])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[216]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[216]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[216]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[216]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[216]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[216]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[216]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[216]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[216].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[217]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [217])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[217]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[217]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[217]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[217]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[217]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[217]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[217]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[217]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[217].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[218]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [218])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[218]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[218]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[218]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[218]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[218]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[218]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[218]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[218]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[218].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[219]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [219])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[219]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[219]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[219]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[219]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[219]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[219]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[219]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[219]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[219].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[220]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [220])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[220]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[220]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[220]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[220]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[220]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[220]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[220]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[220]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[220].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[221]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [221])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[221]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[221]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[221]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[221]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[221]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[221]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[221]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[221]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[221].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[222]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [222])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[222]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[222]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[222]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[222]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[222]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[222]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[222]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[222]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[222].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[223]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [223])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[223]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[223]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[223]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[223]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[223]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[223]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[223]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[223]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[223].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[224]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [224])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[224]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[224]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[224]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[224]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[224]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[224]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[224]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[224]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[224].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[225]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [225])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[225]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[225]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[225]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[225]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[225]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[225]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[225]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[225]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[225].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[226]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [226])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[226]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[226]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[226]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[226]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[226]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[226]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[226]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[226]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[226].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[227]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [227])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[227]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[227]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[227]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[227]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[227]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[227]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[227]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[227]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[227].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[228]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [228])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[228]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[228]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[228]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[228]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[228]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[228]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[228]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[228]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[228].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[229]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [229])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[229]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[229]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[229]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[229]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[229]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[229]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[229]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[229]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[229].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[230]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [230])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[230]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[230]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[230]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[230]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[230]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[230]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[230]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[230]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[230].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[231]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [231])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[231]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[231]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[231]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[231]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[231]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[231]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[231]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[231]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[231].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[232]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [232])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[232]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[232]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[232]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[232]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[232]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[232]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[232]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[232]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[232].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[233]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [233])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[233]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[233]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[233]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[233]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[233]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[233]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[233]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[233]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[233].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[234]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [234])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[234]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[234]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[234]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[234]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[234]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[234]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[234]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[234]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[234].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[235]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [235])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[235]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[235]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[235]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[235]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[235]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[235]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[235]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[235]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[235].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[236]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [236])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[236]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[236]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[236]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[236]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[236]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[236]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[236]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[236]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[236].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[237]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [237])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[237]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[237]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[237]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[237]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[237]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[237]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[237]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[237]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[237].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[238]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [238])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[238]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[238]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[238]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[238]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[238]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[238]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[238]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[238]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[238].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[239]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [239])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[239]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[239]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[239]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[239]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[239]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[239]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[239]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[239]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[239].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[240]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [240])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[240]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[240]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[240]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[240]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[240]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[240]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[240]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[240]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[240].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[241]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [241])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[241]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[241]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[241]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[241]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[241]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[241]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[241]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[241]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[241].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[242]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [242])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[242]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[242]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[242]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[242]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[242]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[242]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[242]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[242]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[242].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[243]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [243])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[243]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[243]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[243]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[243]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[243]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[243]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[243]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[243]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[243].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[244]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [244])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[244]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[244]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[244]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[244]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[244]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[244]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[244]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[244]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[244].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[245]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [245])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[245]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[245]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[245]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[245]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[245]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[245]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[245]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[245]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[245].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[246]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [246])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[246]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[246]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[246]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[246]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[246]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[246]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[246]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[246]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[246].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[247]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [247])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[247]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[247]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[247]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[247]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[247]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[247]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[247]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[247]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[247].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[248]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [248])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[248]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[248]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[248]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[248]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[248]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[248]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[248]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[248]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[248].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[249]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [249])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[249]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[249]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[249]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[249]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[249]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[249]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[249]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[249]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[249].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[250]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [250])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[250]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[250]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[250]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[250]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[250]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[250]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[250]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[250]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[250].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[251]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [251])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[251]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[251]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[251]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[251]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[251]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[251]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[251]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[251]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[251].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[252]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [252])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[252]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[252]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[252]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[252]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[252]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[252]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[252]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[252]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[252].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[253]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [253])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[253]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[253]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[253]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[253]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[253]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[253]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[253]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[253]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[253].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[254]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [254])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[254]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[254]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[254]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[254]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[254]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[254]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[254]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[254]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[254].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[255]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [255])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[255]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[255]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[255]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[255]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[255]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[255]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[255]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clka~FF  (.D(o_pllBr0_reg[255]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[255].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[256]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [256])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[256]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[256]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[256]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[256]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[256]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[256]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[256]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[0]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[256].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[257]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [257])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[257]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[257]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[257]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[257]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[257]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[257]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[257]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[1]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[257].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[258]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [258])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[258]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[258]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[258]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[258]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[258]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[258]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[258]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[2]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[258].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[259]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [259])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[259]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[259]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[259]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[259]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[259]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[259]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[259]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[3]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[259].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[260]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [260])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[260]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[260]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[260]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[260]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[260]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[260]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[260]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[4]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[260].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[261]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [261])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[261]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[261]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[261]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[261]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[261]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[261]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[261]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[5]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[261].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[262]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [262])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[262]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[262]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[262]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[262]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[262]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[262]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[262]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[6]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[262].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[263]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [263])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[263]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[263]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[263]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[263]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[263]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[263]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[263]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[7]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[263].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[264]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [264])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[264]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[264]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[264]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[264]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[264]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[264]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[264]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[8]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[264].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[265]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [265])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[265]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[265]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[265]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[265]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[265]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[265]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[265]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[9]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[265].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[266]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [266])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[266]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[266]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[266]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[266]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[266]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[266]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[266]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[10]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[266].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[267]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [267])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[267]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[267]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[267]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[267]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[267]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[267]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[267]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[11]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[267].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[268]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [268])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[268]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[268]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[268]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[268]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[268]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[268]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[268]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[12]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[268].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[269]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [269])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[269]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[269]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[269]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[269]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[269]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[269]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[269]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[13]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[269].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[270]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [270])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[270]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[270]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[270]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[270]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[270]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[270]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[270]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[14]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[270].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[271]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [271])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[271]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[271]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[271]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[271]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[271]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[271]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[271]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[15]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[271].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[272]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [272])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[272]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[272]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[272]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[272]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[272]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[272]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[272]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[16]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[272].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[273]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [273])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[273]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[273]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[273]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[273]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[273]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[273]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[273]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[17]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[273].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[274]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [274])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[274]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[274]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[274]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[274]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[274]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[274]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[274]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[18]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[274].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[275]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [275])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[275]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[275]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[275]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[275]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[275]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[275]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[275]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[19]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[275].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[276]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [276])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[276]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[276]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[276]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[276]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[276]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[276]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[276]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[20]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[276].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[277]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [277])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[277]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[277]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[277]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[277]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[277]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[277]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[277]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[21]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[277].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[278]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [278])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[278]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[278]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[278]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[278]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[278]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[278]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[278]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[22]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[278].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[279]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [279])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[279]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[279]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[279]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[279]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[279]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[279]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[279]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[23]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[279].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[280]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [280])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[280]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[280]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[280]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[280]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[280]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[280]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[280]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[24]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[280].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[281]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [281])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[281]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[281]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[281]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[281]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[281]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[281]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[281]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[25]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[281].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[282]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [282])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[282]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[282]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[282]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[282]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[282]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[282]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[282]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[26]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[282].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[283]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [283])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[283]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[283]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[283]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[283]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[283]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[283]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[283]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[27]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[283].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[284]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [284])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[284]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[284]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[284]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[284]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[284]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[284]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[284]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[28]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[284].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[285]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [285])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[285]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[285]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[285]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[285]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[285]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[285]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[285]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[29]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[285].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[286]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [286])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[286]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[286]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[286]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[286]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[286]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[286]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[286]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[30]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[286].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[287]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [287])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[287]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[287]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[287]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[287]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[287]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[287]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[287]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[31]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[287].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[288]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [288])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[288]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[288]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[288]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[288]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[288]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[288]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[288]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[32]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[288].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[289]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [289])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[289]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[289]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[289]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[289]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[289]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[289]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[289]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[33]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[289].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[290]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [290])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[290]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[290]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[290]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[290]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[290]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[290]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[290]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[34]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[290].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[291]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [291])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[291]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[291]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[291]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[291]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[291]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[291]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[291]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[35]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[291].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[292]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [292])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[292]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[292]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[292]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[292]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[292]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[292]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[292]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[36]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[292].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[293]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [293])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[293]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[293]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[293]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[293]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[293]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[293]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[293]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[37]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[293].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[294]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [294])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[294]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[294]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[294]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[294]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[294]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[294]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[294]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[38]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[294].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[295]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [295])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[295]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[295]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[295]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[295]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[295]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[295]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[295]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[39]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[295].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[296]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [296])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[296]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[296]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[296]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[296]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[296]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[296]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[296]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[40]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[296].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[297]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [297])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[297]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[297]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[297]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[297]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[297]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[297]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[297]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[41]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[297].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[298]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [298])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[298]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[298]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[298]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[298]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[298]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[298]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[298]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[42]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[298].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[299]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [299])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[299]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[299]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[299]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[299]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[299]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[299]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[299]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[43]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[299].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[300]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [300])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[300]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[300]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[300]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[300]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[300]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[300]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[300]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[44]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[300].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[301]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [301])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[301]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[301]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[301]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[301]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[301]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[301]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[301]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[45]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[301].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[302]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [302])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[302]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[302]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[302]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[302]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[302]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[302]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[302]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[46]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[302].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[303]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [303])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[303]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[303]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[303]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[303]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[303]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[303]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[303]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[47]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[303].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[304]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [304])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[304]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[304]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[304]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[304]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[304]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[304]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[304]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[48]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[304].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[305]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [305])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[305]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[305]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[305]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[305]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[305]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[305]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[305]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[49]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[305].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[306]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [306])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[306]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[306]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[306]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[306]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[306]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[306]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[306]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[50]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[306].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[307]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [307])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[307]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[307]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[307]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[307]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[307]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[307]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[307]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[51]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[307].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[308]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [308])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[308]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[308]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[308]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[308]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[308]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[308]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[308]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[52]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[308].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[309]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [309])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[309]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[309]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[309]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[309]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[309]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[309]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[309]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[53]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[309].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[310]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [310])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[310]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[310]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[310]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[310]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[310]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[310]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[310]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[54]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[310].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[311]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [311])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[311]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[311]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[311]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[311]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[311]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[311]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[311]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[55]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[311].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[312]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [312])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[312]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[312]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[312]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[312]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[312]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[312]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[312]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[56]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[312].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[313]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [313])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[313]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[313]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[313]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[313]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[313]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[313]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[313]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[57]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[313].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[314]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [314])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[314]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[314]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[314]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[314]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[314]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[314]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[314]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[58]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[314].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[315]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [315])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[315]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[315]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[315]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[315]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[315]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[315]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[315]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[59]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[315].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[316]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [316])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[316]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[316]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[316]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[316]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[316]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[316]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[316]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[60]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[316].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[317]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [317])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[317]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[317]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[317]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[317]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[317]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[317]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[317]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[61]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[317].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[318]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [318])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[318]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[318]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[318]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[318]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[318]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[318]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[318]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[62]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[318].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[319]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [319])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[319]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[319]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[319]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[319]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[319]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[319]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[319]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[63]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[319].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[320]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [320])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[320]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[320]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[320]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[320]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[320]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[320]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[320]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[64]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[320].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[321]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [321])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[321]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[321]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[321]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[321]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[321]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[321]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[321]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[65]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[321].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[322]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [322])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[322]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[322]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[322]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[322]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[322]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[322]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[322]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[66]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[322].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[323]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [323])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[323]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[323]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[323]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[323]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[323]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[323]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[323]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[67]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[323].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[324]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [324])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[324]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[324]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[324]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[324]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[324]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[324]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[324]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[68]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[324].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[325]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [325])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[325]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[325]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[325]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[325]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[325]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[325]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[325]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[69]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[325].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[326]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [326])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[326]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[326]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[326]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[326]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[326]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[326]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[326]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[70]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[326].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[327]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [327])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[327]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[327]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[327]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[327]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[327]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[327]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[327]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[71]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[327].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[328]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [328])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[328]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[328]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[328]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[328]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[328]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[328]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[328]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[72]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[328].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[329]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [329])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[329]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[329]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[329]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[329]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[329]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[329]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[329]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[73]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[329].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[330]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [330])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[330]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[330]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[330]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[330]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[330]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[330]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[330]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[74]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[330].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[331]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [331])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[331]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[331]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[331]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[331]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[331]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[331]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[331]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[75]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[331].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[332]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [332])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[332]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[332]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[332]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[332]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[332]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[332]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[332]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[76]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[332].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[333]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [333])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[333]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[333]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[333]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[333]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[333]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[333]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[333]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[77]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[333].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[334]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [334])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[334]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[334]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[334]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[334]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[334]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[334]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[334]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[78]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[334].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[335]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [335])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[335]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[335]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[335]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[335]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[335]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[335]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[335]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[79]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[335].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[336]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [336])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[336]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[336]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[336]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[336]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[336]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[336]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[336]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[80]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[336].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[337]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [337])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[337]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[337]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[337]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[337]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[337]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[337]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[337]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[81]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[337].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[338]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [338])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[338]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[338]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[338]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[338]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[338]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[338]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[338]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[82]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[338].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[339]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [339])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[339]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[339]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[339]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[339]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[339]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[339]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[339]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[83]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[339].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[340]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [340])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[340]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[340]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[340]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[340]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[340]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[340]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[340]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[84]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[340].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[341]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [341])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[341]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[341]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[341]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[341]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[341]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[341]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[341]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[85]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[341].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[342]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [342])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[342]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[342]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[342]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[342]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[342]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[342]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[342]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[86]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[342].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[343]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [343])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[343]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[343]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[343]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[343]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[343]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[343]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[343]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[87]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[343].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[344]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [344])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[344]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[344]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[344]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[344]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[344]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[344]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[344]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[88]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[344].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[345]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [345])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[345]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[345]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[345]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[345]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[345]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[345]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[345]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[89]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[345].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[346]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [346])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[346]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[346]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[346]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[346]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[346]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[346]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[346]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[90]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[346].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[347]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [347])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[347]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[347]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[347]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[347]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[347]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[347]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[347]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[91]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[347].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[348]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [348])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[348]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[348]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[348]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[348]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[348]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[348]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[348]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[92]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[348].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[349]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [349])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[349]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[349]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[349]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[349]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[349]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[349]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[349]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[93]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[349].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[350]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [350])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[350]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[350]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[350]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[350]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[350]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[350]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[350]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[94]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[350].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[351]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [351])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[351]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[351]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[351]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[351]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[351]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[351]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[351]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[95]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[351].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[352]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [352])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[352]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[352]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[352]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[352]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[352]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[352]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[352]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[96]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[352].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[353]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [353])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[353]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[353]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[353]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[353]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[353]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[353]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[353]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[97]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[353].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[354]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [354])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[354]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[354]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[354]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[354]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[354]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[354]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[354]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[98]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[354].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[355]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [355])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[355]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[355]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[355]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[355]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[355]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[355]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[355]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[99]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[355].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[356]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [356])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[356]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[356]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[356]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[356]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[356]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[356]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[356]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[100]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[356].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[357]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [357])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[357]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[357]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[357]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[357]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[357]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[357]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[357]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[101]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[357].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[358]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [358])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[358]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[358]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[358]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[358]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[358]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[358]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[358]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[102]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[358].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[359]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [359])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[359]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[359]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[359]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[359]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[359]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[359]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[359]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[103]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[359].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[360]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [360])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[360]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[360]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[360]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[360]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[360]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[360]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[360]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[104]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[360].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[361]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [361])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[361]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[361]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[361]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[361]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[361]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[361]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[361]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[105]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[361].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[362]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [362])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[362]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[362]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[362]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[362]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[362]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[362]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[362]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[106]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[362].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[363]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [363])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[363]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[363]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[363]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[363]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[363]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[363]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[363]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[107]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[363].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[364]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [364])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[364]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[364]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[364]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[364]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[364]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[364]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[364]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[108]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[364].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[365]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [365])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[365]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[365]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[365]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[365]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[365]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[365]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[365]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[109]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[365].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[366]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [366])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[366]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[366]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[366]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[366]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[366]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[366]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[366]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[110]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[366].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[367]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [367])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[367]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[367]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[367]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[367]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[367]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[367]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[367]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[111]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[367].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[368]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [368])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[368]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[368]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[368]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[368]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[368]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[368]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[368]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[112]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[368].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[369]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [369])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[369]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[369]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[369]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[369]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[369]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[369]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[369]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[113]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[369].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[370]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [370])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[370]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[370]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[370]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[370]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[370]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[370]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[370]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[114]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[370].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[371]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [371])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[371]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[371]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[371]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[371]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[371]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[371]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[371]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[115]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[371].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[372]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [372])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[372]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[372]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[372]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[372]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[372]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[372]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[372]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[116]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[372].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[373]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [373])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[373]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[373]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[373]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[373]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[373]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[373]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[373]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[117]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[373].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[374]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [374])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[374]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[374]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[374]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[374]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[374]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[374]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[374]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[118]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[374].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[375]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [375])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[375]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[375]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[375]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[375]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[375]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[375]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[375]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[119]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[375].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[376]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [376])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[376]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[376]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[376]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[376]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[376]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[376]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[376]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[120]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[376].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[377]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [377])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[377]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[377]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[377]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[377]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[377]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[377]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[377]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[121]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[377].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[378]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [378])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[378]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[378]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[378]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[378]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[378]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[378]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[378]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[122]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[378].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[379]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [379])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[379]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[379]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[379]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[379]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[379]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[379]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[379]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[123]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[379].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[380]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [380])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[380]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[380]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[380]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[380]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[380]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[380]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[380]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[124]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[380].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[381]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [381])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[381]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[381]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[381]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[381]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[381]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[381]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[381]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[125]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[381].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[382]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [382])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[382]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[382]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[382]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[382]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[382]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[382]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[382]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[126]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[382].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[383]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [383])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[383]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[383]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[383]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[383]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[383]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[383]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[383]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[127]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[383].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[384]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [384])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[384]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[384]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[384]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[384]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[384]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[384]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[384]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[128]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[384].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[385]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [385])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[385]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[385]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[385]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[385]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[385]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[385]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[385]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[129]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[385].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[386]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [386])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[386]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[386]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[386]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[386]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[386]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[386]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[386]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[130]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[386].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[387]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [387])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[387]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[387]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[387]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[387]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[387]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[387]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[387]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[131]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[387].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[388]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [388])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[388]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[388]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[388]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[388]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[388]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[388]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[388]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[132]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[388].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[389]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [389])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[389]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[389]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[389]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[389]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[389]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[389]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[389]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[133]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[389].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[390]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [390])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[390]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[390]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[390]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[390]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[390]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[390]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[390]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[134]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[390].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[391]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [391])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[391]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[391]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[391]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[391]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[391]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[391]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[391]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[135]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[391].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[392]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [392])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[392]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[392]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[392]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[392]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[392]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[392]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[392]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[136]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[392].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[393]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [393])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[393]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[393]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[393]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[393]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[393]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[393]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[393]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[137]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[393].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[394]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [394])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[394]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[394]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[394]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[394]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[394]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[394]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[394]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[138]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[394].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[395]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [395])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[395]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[395]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[395]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[395]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[395]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[395]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[395]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[139]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[395].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[396]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [396])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[396]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[396]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[396]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[396]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[396]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[396]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[396]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[140]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[396].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[397]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [397])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[397]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[397]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[397]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[397]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[397]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[397]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[397]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[141]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[397].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[398]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [398])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[398]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[398]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[398]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[398]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[398]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[398]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[398]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[142]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[398].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[399]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [399])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[399]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[399]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[399]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[399]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[399]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[399]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[399]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[143]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[399].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[400]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [400])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[400]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[400]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[400]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[400]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[400]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[400]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[400]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[144]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[400].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[401]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [401])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[401]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[401]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[401]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[401]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[401]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[401]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[401]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[145]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[401].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[402]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [402])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[402]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[402]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[402]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[402]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[402]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[402]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[402]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[146]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[402].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[403]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [403])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[403]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[403]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[403]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[403]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[403]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[403]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[403]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[147]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[403].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[404]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [404])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[404]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[404]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[404]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[404]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[404]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[404]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[404]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[148]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[404].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[405]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [405])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[405]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[405]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[405]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[405]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[405]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[405]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[405]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[149]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[405].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[406]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [406])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[406]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[406]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[406]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[406]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[406]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[406]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[406]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[150]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[406].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[407]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [407])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[407]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[407]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[407]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[407]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[407]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[407]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[407]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[151]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[407].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[408]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [408])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[408]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[408]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[408]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[408]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[408]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[408]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[408]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[152]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[408].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[409]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [409])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[409]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[409]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[409]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[409]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[409]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[409]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[409]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[153]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[409].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[410]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [410])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[410]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[410]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[410]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[410]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[410]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[410]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[410]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[154]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[410].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[411]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [411])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[411]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[411]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[411]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[411]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[411]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[411]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[411]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[155]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[411].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[412]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [412])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[412]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[412]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[412]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[412]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[412]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[412]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[412]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[156]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[412].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[413]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [413])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[413]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[413]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[413]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[413]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[413]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[413]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[413]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[157]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[413].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[414]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [414])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[414]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[414]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[414]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[414]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[414]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[414]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[414]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[158]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[414].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[415]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [415])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[415]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[415]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[415]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[415]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[415]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[415]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[415]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[159]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[415].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[416]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [416])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[416]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[416]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[416]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[416]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[416]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[416]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[416]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[160]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[416].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[417]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [417])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[417]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[417]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[417]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[417]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[417]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[417]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[417]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[161]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[417].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[418]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [418])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[418]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[418]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[418]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[418]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[418]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[418]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[418]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[162]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[418].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[419]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [419])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[419]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[419]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[419]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[419]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[419]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[419]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[419]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[163]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[419].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[420]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [420])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[420]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[420]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[420]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[420]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[420]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[420]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[420]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[164]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[420].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[421]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [421])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[421]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[421]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[421]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[421]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[421]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[421]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[421]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[165]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[421].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[422]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [422])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[422]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[422]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[422]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[422]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[422]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[422]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[422]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[166]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[422].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[423]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [423])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[423]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[423]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[423]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[423]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[423]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[423]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[423]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[167]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[423].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[424]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [424])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[424]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[424]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[424]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[424]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[424]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[424]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[424]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[168]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[424].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[425]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [425])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[425]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[425]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[425]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[425]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[425]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[425]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[425]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[169]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[425].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[426]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [426])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[426]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[426]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[426]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[426]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[426]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[426]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[426]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[170]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[426].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[427]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [427])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[427]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[427]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[427]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[427]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[427]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[427]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[427]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[171]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[427].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[428]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [428])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[428]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[428]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[428]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[428]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[428]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[428]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[428]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[172]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[428].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[429]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [429])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[429]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[429]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[429]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[429]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[429]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[429]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[429]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[173]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[429].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[430]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [430])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[430]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[430]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[430]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[430]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[430]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[430]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[430]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[174]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[430].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[431]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [431])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[431]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[431]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[431]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[431]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[431]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[431]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[431]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[175]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[431].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[432]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [432])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[432]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[432]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[432]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[432]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[432]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[432]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[432]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[176]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[432].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[433]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [433])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[433]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[433]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[433]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[433]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[433]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[433]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[433]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[177]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[433].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[434]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [434])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[434]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[434]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[434]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[434]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[434]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[434]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[434]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[178]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[434].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[435]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [435])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[435]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[435]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[435]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[435]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[435]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[435]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[435]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[179]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[435].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[436]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [436])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[436]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[436]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[436]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[436]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[436]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[436]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[436]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[180]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[436].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[437]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [437])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[437]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[437]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[437]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[437]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[437]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[437]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[437]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[181]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[437].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[438]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [438])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[438]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[438]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[438]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[438]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[438]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[438]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[438]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[182]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[438].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[439]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [439])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[439]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[439]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[439]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[439]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[439]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[439]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[439]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[183]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[439].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[440]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [440])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[440]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[440]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[440]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[440]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[440]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[440]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[440]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[184]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[440].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[441]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [441])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[441]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[441]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[441]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[441]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[441]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[441]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[441]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[185]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[441].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[442]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [442])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[442]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[442]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[442]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[442]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[442]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[442]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[442]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[186]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[442].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[443]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [443])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[443]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[443]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[443]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[443]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[443]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[443]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[443]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[187]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[443].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[444]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [444])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[444]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[444]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[444]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[444]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[444]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[444]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[444]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[188]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[444].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[445]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [445])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[445]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[445]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[445]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[445]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[445]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[445]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[445]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[189]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[445].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[446]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [446])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[446]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[446]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[446]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[446]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[446]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[446]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[446]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[190]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[446].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[447]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [447])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[447]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[447]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[447]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[447]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[447]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[447]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[447]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[191]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[447].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[448]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [448])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[448]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[448]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[448]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[448]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[448]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[448]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[448]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[192]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[448].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[449]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [449])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[449]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[449]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[449]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[449]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[449]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[449]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[449]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[193]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[449].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[450]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [450])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[450]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[450]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[450]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[450]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[450]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[450]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[450]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[194]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[450].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[451]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [451])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[451]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[451]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[451]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[451]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[451]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[451]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[451]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[195]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[451].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[452]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [452])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[452]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[452]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[452]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[452]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[452]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[452]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[452]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[196]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[452].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[453]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [453])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[453]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[453]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[453]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[453]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[453]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[453]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[453]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[197]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[453].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[454]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [454])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[454]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[454]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[454]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[454]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[454]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[454]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[454]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[198]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[454].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[455]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [455])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[455]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[455]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[455]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[455]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[455]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[455]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[455]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[199]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[455].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[456]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [456])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[456]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[456]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[456]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[456]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[456]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[456]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[456]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[200]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[456].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[457]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [457])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[457]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[457]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[457]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[457]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[457]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[457]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[457]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[201]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[457].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[458]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [458])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[458]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[458]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[458]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[458]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[458]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[458]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[458]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[202]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[458].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[459]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [459])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[459]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[459]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[459]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[459]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[459]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[459]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[459]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[203]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[459].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[460]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [460])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[460]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[460]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[460]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[460]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[460]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[460]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[460]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[204]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[460].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[461]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [461])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[461]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[461]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[461]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[461]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[461]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[461]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[461]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[205]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[461].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[462]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [462])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[462]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[462]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[462]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[462]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[462]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[462]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[462]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[206]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[462].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[463]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [463])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[463]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[463]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[463]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[463]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[463]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[463]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[463]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[207]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[463].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[464]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [464])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[464]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[464]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[464]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[464]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[464]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[464]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[464]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[208]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[464].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[465]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [465])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[465]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[465]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[465]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[465]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[465]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[465]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[465]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[209]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[465].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[466]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [466])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[466]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[466]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[466]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[466]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[466]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[466]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[466]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[210]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[466].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[467]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [467])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[467]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[467]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[467]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[467]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[467]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[467]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[467]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[211]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[467].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[468]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [468])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[468]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[468]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[468]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[468]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[468]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[468]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[468]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[212]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[468].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[469]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [469])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[469]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[469]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[469]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[469]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[469]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[469]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[469]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[213]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[469].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[470]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [470])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[470]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[470]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[470]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[470]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[470]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[470]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[470]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[214]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[470].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[471]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [471])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[471]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[471]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[471]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[471]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[471]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[471]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[471]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[215]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[471].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[472]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [472])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[472]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[472]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[472]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[472]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[472]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[472]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[472]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[216]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[472].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[473]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [473])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[473]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[473]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[473]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[473]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[473]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[473]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[473]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[217]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[473].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[474]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [474])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[474]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[474]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[474]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[474]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[474]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[474]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[474]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[218]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[474].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[475]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [475])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[475]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[475]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[475]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[475]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[475]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[475]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[475]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[219]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[475].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[476]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [476])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[476]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[476]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[476]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[476]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[476]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[476]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[476]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[220]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[476].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[477]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [477])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[477]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[477]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[477]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[477]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[477]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[477]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[477]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[221]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[477].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[478]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [478])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[478]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[478]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[478]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[478]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[478]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[478]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[478]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[222]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[478].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[479]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [479])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[479]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[479]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[479]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[479]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[479]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[479]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[479]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[223]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[479].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[480]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [480])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[480]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[480]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[480]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[480]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[480]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[480]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[480]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[224]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[480].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[481]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [481])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[481]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[481]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[481]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[481]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[481]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[481]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[481]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[225]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[481].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[482]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [482])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[482]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[482]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[482]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[482]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[482]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[482]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[482]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[226]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[482].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[483]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [483])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[483]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[483]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[483]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[483]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[483]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[483]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[483]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[227]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[483].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[484]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [484])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[484]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[484]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[484]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[484]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[484]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[484]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[484]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[228]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[484].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[485]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [485])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[485]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[485]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[485]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[485]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[485]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[485]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[485]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[229]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[485].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[486]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [486])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[486]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[486]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[486]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[486]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[486]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[486]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[486]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[230]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[486].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[487]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [487])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[487]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[487]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[487]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[487]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[487]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[487]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[487]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[231]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[487].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[488]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [488])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[488]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[488]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[488]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[488]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[488]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[488]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[488]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[232]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[488].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[489]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [489])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[489]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[489]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[489]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[489]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[489]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[489]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[489]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[233]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[489].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[490]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [490])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[490]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[490]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[490]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[490]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[490]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[490]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[490]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[234]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[490].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[491]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [491])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[491]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[491]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[491]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[491]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[491]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[491]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[491]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[235]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[491].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[492]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [492])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[492]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[492]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[492]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[492]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[492]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[492]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[492]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[236]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[492].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[493]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [493])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[493]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[493]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[493]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[493]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[493]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[493]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[493]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[237]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[493].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[494]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [494])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[494]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[494]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[494]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[494]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[494]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[494]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[494]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[238]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[494].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[495]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [495])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[495]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[495]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[495]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[495]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[495]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[495]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[495]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[239]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[495].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[496]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [496])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[496]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[496]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[496]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[496]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[496]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[496]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[496]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[240]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[496].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[497]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [497])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[497]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[497]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[497]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[497]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[497]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[497]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[497]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[241]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[497].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[498]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [498])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[498]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[498]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[498]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[498]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[498]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[498]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[498]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[242]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[498].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[499]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [499])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[499]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[499]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[499]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[499]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[499]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[499]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[499]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[243]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[499].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[500]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [500])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[500]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[500]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[500]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[500]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[500]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[500]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[500]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[244]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[500].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[501]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [501])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[501]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[501]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[501]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[501]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[501]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[501]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[501]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[245]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[501].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[502]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [502])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[502]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[502]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[502]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[502]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[502]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[502]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[502]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[246]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[502].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[503]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [503])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[503]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[503]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[503]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[503]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[503]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[503]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[503]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[247]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[503].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[504]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [504])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[504]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[504]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[504]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[504]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[504]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[504]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[504]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[248]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[504].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[505]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [505])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[505]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[505]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[505]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[505]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[505]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[505]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[505]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[249]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[505].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[506]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [506])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[506]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[506]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[506]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[506]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[506]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[506]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[506]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[250]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[506].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[507]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [507])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[507]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[507]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[507]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[507]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[507]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[507]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[507]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[251]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[507].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[508]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [508])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[508]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[508]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[508]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[508]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[508]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[508]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[508]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[252]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[508].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[509]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [509])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[509]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[509]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[509]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[509]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[509]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[509]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[509]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[253]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[509].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[510]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [510])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[510]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[510]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[510]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[510]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[510]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[510]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[510]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[254]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[510].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clkb~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clka ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clkb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clkb~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clkb~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clkb~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clkb~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clkb~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clkb~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clkb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/probe_in_sync[511]~FF  (.D(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clkb ), 
           .CE(1'b1), .CLK(\clk_0~O ), .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/probe_in_sync [511])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1905)
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[511]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[511]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[511]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[511]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[511]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[511]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/probe_in_sync[511]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clka~FF  (.D(o_pllBr1_reg[255]), 
           .CE(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), .CLK(\bscan_TCK~O ), 
           .SR(1'b0), .Q(\debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clka )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1894)
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clka~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clka~FF .CE_POLARITY = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clka~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clka~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clka~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clka~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/gen_probe_in_sync[511].sync_probe_in_U/d_clka~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/internal_register_select[1]~FF  (.D(\debug_inst/edb_user_dr [74]), 
           .CE(\debug_inst/vio0/vio_core_inst/regsel_ld_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/internal_register_select [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1351)
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[1]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[1]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[1]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[1]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[1]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[1]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/internal_register_select[2]~FF  (.D(\debug_inst/edb_user_dr [75]), 
           .CE(\debug_inst/vio0/vio_core_inst/regsel_ld_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/internal_register_select [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1351)
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[2]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[2]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[2]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[2]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[2]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[2]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/vio0/vio_core_inst/internal_register_select[3]~FF  (.D(\debug_inst/edb_user_dr [76]), 
           .CE(\debug_inst/vio0/vio_core_inst/regsel_ld_en ), .CLK(\bscan_TCK~O ), 
           .SR(\debug_inst/edb_soft_reset ), .Q(\debug_inst/vio0/vio_core_inst/internal_register_select [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1351)
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[3]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[3]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[3]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[3]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[3]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[3]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/vio0/vio_core_inst/internal_register_select[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/debug_hub_inst/module_id_reg[0]~FF  (.D(\debug_inst/edb_user_dr [77]), 
           .CE(\debug_inst/debug_hub_inst/n267 ), .CLK(\bscan_TCK~O ), .SR(1'b0), 
           .Q(\debug_inst/debug_hub_inst/module_id_reg [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(437)
    defparam \debug_inst/debug_hub_inst/module_id_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_soft_reset~FF  (.D(\debug_inst/edb_user_dr [76]), 
           .CE(\debug_inst/debug_hub_inst/n265 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_soft_reset )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(443)
    defparam \debug_inst/edb_soft_reset~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_soft_reset~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_soft_reset~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_soft_reset~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_soft_reset~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_soft_reset~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_soft_reset~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/debug_hub_inst/module_id_reg[1]~FF  (.D(\debug_inst/edb_user_dr [78]), 
           .CE(\debug_inst/debug_hub_inst/n267 ), .CLK(\bscan_TCK~O ), .SR(1'b0), 
           .Q(\debug_inst/debug_hub_inst/module_id_reg [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(437)
    defparam \debug_inst/debug_hub_inst/module_id_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/debug_hub_inst/module_id_reg[2]~FF  (.D(\debug_inst/edb_user_dr [79]), 
           .CE(\debug_inst/debug_hub_inst/n267 ), .CLK(\bscan_TCK~O ), .SR(1'b0), 
           .Q(\debug_inst/debug_hub_inst/module_id_reg [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(437)
    defparam \debug_inst/debug_hub_inst/module_id_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/debug_hub_inst/module_id_reg[3]~FF  (.D(\debug_inst/edb_user_dr [80]), 
           .CE(\debug_inst/debug_hub_inst/n267 ), .CLK(\bscan_TCK~O ), .SR(1'b0), 
           .Q(\debug_inst/debug_hub_inst/module_id_reg [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(437)
    defparam \debug_inst/debug_hub_inst/module_id_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC = 1'b1;
    defparam \debug_inst/debug_hub_inst/module_id_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[45]~FF  (.D(\debug_inst/edb_user_dr [46]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[45]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[45]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[45]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[45]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[45]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[45]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[46]~FF  (.D(\debug_inst/edb_user_dr [47]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[46]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[46]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[46]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[46]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[46]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[46]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[47]~FF  (.D(\debug_inst/edb_user_dr [48]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[47]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[47]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[47]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[47]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[47]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[47]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[48]~FF  (.D(\debug_inst/edb_user_dr [49]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[48]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[48]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[48]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[48]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[48]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[48]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[49]~FF  (.D(\debug_inst/edb_user_dr [50]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[49]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[49]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[49]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[49]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[49]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[49]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[50]~FF  (.D(\debug_inst/edb_user_dr [51]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[50]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[50]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[50]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[50]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[50]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[50]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[51]~FF  (.D(\debug_inst/edb_user_dr [52]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[51]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[51]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[51]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[51]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[51]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[51]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[52]~FF  (.D(\debug_inst/edb_user_dr [53]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[52]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[52]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[52]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[52]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[52]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[52]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[53]~FF  (.D(\debug_inst/edb_user_dr [54]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[53]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[53]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[53]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[53]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[53]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[53]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[54]~FF  (.D(\debug_inst/edb_user_dr [55]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[54]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[54]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[54]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[54]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[54]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[54]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[55]~FF  (.D(\debug_inst/edb_user_dr [56]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[55]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[55]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[55]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[55]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[55]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[55]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[56]~FF  (.D(\debug_inst/edb_user_dr [57]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[56]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[56]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[56]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[56]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[56]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[56]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[57]~FF  (.D(\debug_inst/edb_user_dr [58]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[57]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[57]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[57]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[57]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[57]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[57]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[58]~FF  (.D(\debug_inst/edb_user_dr [59]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[58]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[58]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[58]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[58]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[58]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[58]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[59]~FF  (.D(\debug_inst/edb_user_dr [60]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[59]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[59]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[59]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[59]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[59]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[59]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[60]~FF  (.D(\debug_inst/edb_user_dr [61]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [60])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[60]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[60]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[60]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[60]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[60]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[60]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[61]~FF  (.D(\debug_inst/edb_user_dr [62]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [61])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[61]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[61]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[61]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[61]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[61]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[61]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[62]~FF  (.D(\debug_inst/edb_user_dr [63]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [62])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[62]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[62]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[62]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[62]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[62]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[62]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[63]~FF  (.D(\debug_inst/edb_user_dr [64]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [63])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[63]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[63]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[63]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[63]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[63]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[63]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[64]~FF  (.D(\debug_inst/edb_user_dr [65]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [64])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[64]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[64]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[64]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[64]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[64]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[64]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[65]~FF  (.D(\debug_inst/edb_user_dr [66]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [65])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[65]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[65]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[65]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[65]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[65]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[65]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[66]~FF  (.D(\debug_inst/edb_user_dr [67]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [66])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[66]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[66]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[66]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[66]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[66]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[66]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[67]~FF  (.D(\debug_inst/edb_user_dr [68]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [67])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[67]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[67]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[67]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[67]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[67]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[67]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[68]~FF  (.D(\debug_inst/edb_user_dr [69]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [68])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[68]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[68]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[68]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[68]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[68]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[68]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[69]~FF  (.D(\debug_inst/edb_user_dr [70]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [69])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[69]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[69]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[69]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[69]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[69]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[69]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[70]~FF  (.D(\debug_inst/edb_user_dr [71]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [70])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[70]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[70]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[70]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[70]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[70]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[70]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[71]~FF  (.D(\debug_inst/edb_user_dr [72]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [71])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[71]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[71]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[71]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[71]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[71]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[71]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[72]~FF  (.D(\debug_inst/edb_user_dr [73]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [72])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[72]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[72]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[72]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[72]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[72]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[72]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[73]~FF  (.D(\debug_inst/edb_user_dr [74]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [73])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[73]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[73]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[73]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[73]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[73]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[73]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[74]~FF  (.D(\debug_inst/edb_user_dr [75]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [74])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[74]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[74]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[74]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[74]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[74]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[74]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[75]~FF  (.D(\debug_inst/edb_user_dr [76]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [75])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[75]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[75]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[75]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[75]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[75]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[75]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[76]~FF  (.D(\debug_inst/edb_user_dr [77]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [76])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[76]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[76]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[76]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[76]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[76]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[76]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[77]~FF  (.D(\debug_inst/edb_user_dr [78]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [77])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[77]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[77]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[77]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[77]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[77]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[77]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[78]~FF  (.D(\debug_inst/edb_user_dr [79]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [78])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[78]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[78]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[78]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[78]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[78]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[78]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[79]~FF  (.D(\debug_inst/edb_user_dr [80]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [79])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[79]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[79]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[79]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[79]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[79]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[79]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[80]~FF  (.D(\debug_inst/edb_user_dr [81]), 
           .CE(\debug_inst/debug_hub_inst/n96 ), .CLK(\bscan_TCK~O ), .SR(bscan_RESET), 
           .Q(\debug_inst/edb_user_dr [80])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[80]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[80]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[80]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[80]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[80]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[80]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \debug_inst/edb_user_dr[81]~FF  (.D(bscan_TDI), .CE(\debug_inst/debug_hub_inst/n96 ), 
           .CLK(\bscan_TCK~O ), .SR(bscan_RESET), .Q(\debug_inst/edb_user_dr [81])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(429)
    defparam \debug_inst/edb_user_dr[81]~FF .CLK_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[81]~FF .CE_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[81]~FF .SR_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[81]~FF .D_POLARITY = 1'b1;
    defparam \debug_inst/edb_user_dr[81]~FF .SR_SYNC = 1'b0;
    defparam \debug_inst/edb_user_dr[81]~FF .SR_VALUE = 1'b0;
    defparam \debug_inst/edb_user_dr[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \test_module/add_41/i90  (.I0(o_pllBr0_reg[90]), .I1(1'b0), 
            .CI(\test_module/add_41/n178 ), .O(\test_module/n33 [90]), .CO(\test_module/add_41/n180 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i90 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i90 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i86  (.I0(o_pllBr0_reg[86]), .I1(1'b0), 
            .CI(\test_module/add_41/n170 ), .O(\test_module/n33 [86]), .CO(\test_module/add_41/n172 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i86 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i86 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i95  (.I0(o_pllBr0_reg[95]), .I1(1'b0), 
            .CI(\test_module/add_41/n188 ), .O(\test_module/n33 [95]), .CO(\test_module/add_41/n190 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i95 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i95 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i1  (.I0(o_pllBr0_reg[1]), .I1(o_pllBr0_reg[0]), 
            .CI(1'b0), .O(\test_module/n33 [1]), .CO(\test_module/add_41/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i1 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i85  (.I0(o_pllBr0_reg[85]), .I1(1'b0), 
            .CI(\test_module/add_41/n168 ), .O(\test_module/n33 [85]), .CO(\test_module/add_41/n170 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i85 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i85 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_44/i1  (.I0(\test_module/delay_2 [1]), .I1(\test_module/delay_2 [0]), 
            .CI(1'b0), .O(\test_module/n1132 [1]), .CO(\test_module/add_44/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(34)
    defparam \test_module/add_44/i1 .I0_POLARITY = 1'b1;
    defparam \test_module/add_44/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i96  (.I0(o_pllBr0_reg[96]), .I1(1'b0), 
            .CI(\test_module/add_41/n190 ), .O(\test_module/n33 [96]), .CO(\test_module/add_41/n192 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i96 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i96 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i84  (.I0(o_pllBr0_reg[84]), .I1(1'b0), 
            .CI(\test_module/add_41/n166 ), .O(\test_module/n33 [84]), .CO(\test_module/add_41/n168 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i84 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i84 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i83  (.I0(o_pllBr0_reg[83]), .I1(1'b0), 
            .CI(\test_module/add_41/n164 ), .O(\test_module/n33 [83]), .CO(\test_module/add_41/n166 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i83 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i83 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i1  (.I0(o_pllBr1_reg[1]), .I1(o_pllBr1_reg[0]), 
            .CI(1'b0), .O(\test_module/n1156 [1]), .CO(\test_module/add_46/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i1 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \debug_inst/vio0/vio_core_inst/add_772/i1  (.I0(\debug_inst/vio0/vio_core_inst/bit_count [1]), 
            .I1(\debug_inst/vio0/vio_core_inst/bit_count [0]), .CI(1'b0), 
            .O(\debug_inst/vio0/vio_core_inst/n408 [1]), .CO(\debug_inst/vio0/vio_core_inst/add_772/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1429)
    defparam \debug_inst/vio0/vio_core_inst/add_772/i1 .I0_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/add_772/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i97  (.I0(o_pllBr0_reg[97]), .I1(1'b0), 
            .CI(\test_module/add_41/n192 ), .O(\test_module/n33 [97]), .CO(\test_module/add_41/n194 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i97 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i97 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i82  (.I0(o_pllBr0_reg[82]), .I1(1'b0), 
            .CI(\test_module/add_41/n162 ), .O(\test_module/n33 [82]), .CO(\test_module/add_41/n164 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i82 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i82 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i81  (.I0(o_pllBr0_reg[81]), .I1(1'b0), 
            .CI(\test_module/add_41/n160 ), .O(\test_module/n33 [81]), .CO(\test_module/add_41/n162 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i81 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i81 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i80  (.I0(o_pllBr0_reg[80]), .I1(1'b0), 
            .CI(\test_module/add_41/n158 ), .O(\test_module/n33 [80]), .CO(\test_module/add_41/n160 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i80 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i80 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i79  (.I0(o_pllBr0_reg[79]), .I1(1'b0), 
            .CI(\test_module/add_41/n156 ), .O(\test_module/n33 [79]), .CO(\test_module/add_41/n158 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i79 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i79 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i78  (.I0(o_pllBr0_reg[78]), .I1(1'b0), 
            .CI(\test_module/add_41/n154 ), .O(\test_module/n33 [78]), .CO(\test_module/add_41/n156 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i78 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i78 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i77  (.I0(o_pllBr0_reg[77]), .I1(1'b0), 
            .CI(\test_module/add_41/n152 ), .O(\test_module/n33 [77]), .CO(\test_module/add_41/n154 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i77 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i77 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i76  (.I0(o_pllBr0_reg[76]), .I1(1'b0), 
            .CI(\test_module/add_41/n150 ), .O(\test_module/n33 [76]), .CO(\test_module/add_41/n152 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i76 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i76 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i75  (.I0(o_pllBr0_reg[75]), .I1(1'b0), 
            .CI(\test_module/add_41/n148 ), .O(\test_module/n33 [75]), .CO(\test_module/add_41/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i75 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i75 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i74  (.I0(o_pllBr0_reg[74]), .I1(1'b0), 
            .CI(\test_module/add_41/n146 ), .O(\test_module/n33 [74]), .CO(\test_module/add_41/n148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i74 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i74 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i98  (.I0(o_pllBr0_reg[98]), .I1(1'b0), 
            .CI(\test_module/add_41/n194 ), .O(\test_module/n33 [98]), .CO(\test_module/add_41/n196 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i98 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i98 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i99  (.I0(o_pllBr0_reg[99]), .I1(1'b0), 
            .CI(\test_module/add_41/n196 ), .O(\test_module/n33 [99]), .CO(\test_module/add_41/n198 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i99 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i99 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i100  (.I0(o_pllBr0_reg[100]), .I1(1'b0), 
            .CI(\test_module/add_41/n198 ), .O(\test_module/n33 [100]), 
            .CO(\test_module/add_41/n200 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i100 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i100 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i101  (.I0(o_pllBr0_reg[101]), .I1(1'b0), 
            .CI(\test_module/add_41/n200 ), .O(\test_module/n33 [101]), 
            .CO(\test_module/add_41/n202 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i101 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i101 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i102  (.I0(o_pllBr0_reg[102]), .I1(1'b0), 
            .CI(\test_module/add_41/n202 ), .O(\test_module/n33 [102]), 
            .CO(\test_module/add_41/n204 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i102 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i102 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i103  (.I0(o_pllBr0_reg[103]), .I1(1'b0), 
            .CI(\test_module/add_41/n204 ), .O(\test_module/n33 [103]), 
            .CO(\test_module/add_41/n206 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i103 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i103 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i104  (.I0(o_pllBr0_reg[104]), .I1(1'b0), 
            .CI(\test_module/add_41/n206 ), .O(\test_module/n33 [104]), 
            .CO(\test_module/add_41/n208 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i104 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i104 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i105  (.I0(o_pllBr0_reg[105]), .I1(1'b0), 
            .CI(\test_module/add_41/n208 ), .O(\test_module/n33 [105]), 
            .CO(\test_module/add_41/n210 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i105 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i105 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i106  (.I0(o_pllBr0_reg[106]), .I1(1'b0), 
            .CI(\test_module/add_41/n210 ), .O(\test_module/n33 [106]), 
            .CO(\test_module/add_41/n212 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i106 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i106 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i107  (.I0(o_pllBr0_reg[107]), .I1(1'b0), 
            .CI(\test_module/add_41/n212 ), .O(\test_module/n33 [107]), 
            .CO(\test_module/add_41/n214 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i107 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i107 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i108  (.I0(o_pllBr0_reg[108]), .I1(1'b0), 
            .CI(\test_module/add_41/n214 ), .O(\test_module/n33 [108]), 
            .CO(\test_module/add_41/n216 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i108 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i108 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i109  (.I0(o_pllBr0_reg[109]), .I1(1'b0), 
            .CI(\test_module/add_41/n216 ), .O(\test_module/n33 [109]), 
            .CO(\test_module/add_41/n218 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i109 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i109 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i110  (.I0(o_pllBr0_reg[110]), .I1(1'b0), 
            .CI(\test_module/add_41/n218 ), .O(\test_module/n33 [110]), 
            .CO(\test_module/add_41/n220 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i110 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i110 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i111  (.I0(o_pllBr0_reg[111]), .I1(1'b0), 
            .CI(\test_module/add_41/n220 ), .O(\test_module/n33 [111]), 
            .CO(\test_module/add_41/n222 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i111 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i111 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i112  (.I0(o_pllBr0_reg[112]), .I1(1'b0), 
            .CI(\test_module/add_41/n222 ), .O(\test_module/n33 [112]), 
            .CO(\test_module/add_41/n224 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i112 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i112 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i113  (.I0(o_pllBr0_reg[113]), .I1(1'b0), 
            .CI(\test_module/add_41/n224 ), .O(\test_module/n33 [113]), 
            .CO(\test_module/add_41/n226 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i113 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i113 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i114  (.I0(o_pllBr0_reg[114]), .I1(1'b0), 
            .CI(\test_module/add_41/n226 ), .O(\test_module/n33 [114]), 
            .CO(\test_module/add_41/n228 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i114 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i114 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i115  (.I0(o_pllBr0_reg[115]), .I1(1'b0), 
            .CI(\test_module/add_41/n228 ), .O(\test_module/n33 [115]), 
            .CO(\test_module/add_41/n230 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i115 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i115 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i116  (.I0(o_pllBr0_reg[116]), .I1(1'b0), 
            .CI(\test_module/add_41/n230 ), .O(\test_module/n33 [116]), 
            .CO(\test_module/add_41/n232 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i116 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i116 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i117  (.I0(o_pllBr0_reg[117]), .I1(1'b0), 
            .CI(\test_module/add_41/n232 ), .O(\test_module/n33 [117]), 
            .CO(\test_module/add_41/n234 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i117 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i117 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i118  (.I0(o_pllBr0_reg[118]), .I1(1'b0), 
            .CI(\test_module/add_41/n234 ), .O(\test_module/n33 [118]), 
            .CO(\test_module/add_41/n236 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i118 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i118 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i73  (.I0(o_pllBr0_reg[73]), .I1(1'b0), 
            .CI(\test_module/add_41/n144 ), .O(\test_module/n33 [73]), .CO(\test_module/add_41/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i73 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i73 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i72  (.I0(o_pllBr0_reg[72]), .I1(1'b0), 
            .CI(\test_module/add_41/n142 ), .O(\test_module/n33 [72]), .CO(\test_module/add_41/n144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i72 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i72 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i71  (.I0(o_pllBr0_reg[71]), .I1(1'b0), 
            .CI(\test_module/add_41/n140 ), .O(\test_module/n33 [71]), .CO(\test_module/add_41/n142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i71 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i71 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i70  (.I0(o_pllBr0_reg[70]), .I1(1'b0), 
            .CI(\test_module/add_41/n138 ), .O(\test_module/n33 [70]), .CO(\test_module/add_41/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i70 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i70 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i69  (.I0(o_pllBr0_reg[69]), .I1(1'b0), 
            .CI(\test_module/add_41/n136 ), .O(\test_module/n33 [69]), .CO(\test_module/add_41/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i69 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i69 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i68  (.I0(o_pllBr0_reg[68]), .I1(1'b0), 
            .CI(\test_module/add_41/n134 ), .O(\test_module/n33 [68]), .CO(\test_module/add_41/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i68 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i68 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i67  (.I0(o_pllBr0_reg[67]), .I1(1'b0), 
            .CI(\test_module/add_41/n132 ), .O(\test_module/n33 [67]), .CO(\test_module/add_41/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i67 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i67 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i119  (.I0(o_pllBr0_reg[119]), .I1(1'b0), 
            .CI(\test_module/add_41/n236 ), .O(\test_module/n33 [119]), 
            .CO(\test_module/add_41/n238 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i119 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i119 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i120  (.I0(o_pllBr0_reg[120]), .I1(1'b0), 
            .CI(\test_module/add_41/n238 ), .O(\test_module/n33 [120]), 
            .CO(\test_module/add_41/n240 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i120 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i120 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i121  (.I0(o_pllBr0_reg[121]), .I1(1'b0), 
            .CI(\test_module/add_41/n240 ), .O(\test_module/n33 [121]), 
            .CO(\test_module/add_41/n242 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i121 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i121 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i122  (.I0(o_pllBr0_reg[122]), .I1(1'b0), 
            .CI(\test_module/add_41/n242 ), .O(\test_module/n33 [122]), 
            .CO(\test_module/add_41/n244 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i122 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i122 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i123  (.I0(o_pllBr0_reg[123]), .I1(1'b0), 
            .CI(\test_module/add_41/n244 ), .O(\test_module/n33 [123]), 
            .CO(\test_module/add_41/n246 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i123 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i123 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i124  (.I0(o_pllBr0_reg[124]), .I1(1'b0), 
            .CI(\test_module/add_41/n246 ), .O(\test_module/n33 [124]), 
            .CO(\test_module/add_41/n248 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i124 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i124 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i125  (.I0(o_pllBr0_reg[125]), .I1(1'b0), 
            .CI(\test_module/add_41/n248 ), .O(\test_module/n33 [125]), 
            .CO(\test_module/add_41/n250 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i125 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i125 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i126  (.I0(o_pllBr0_reg[126]), .I1(1'b0), 
            .CI(\test_module/add_41/n250 ), .O(\test_module/n33 [126]), 
            .CO(\test_module/add_41/n252 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i126 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i126 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i127  (.I0(o_pllBr0_reg[127]), .I1(1'b0), 
            .CI(\test_module/add_41/n252 ), .O(\test_module/n33 [127]), 
            .CO(\test_module/add_41/n254 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i127 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i127 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i128  (.I0(o_pllBr0_reg[128]), .I1(1'b0), 
            .CI(\test_module/add_41/n254 ), .O(\test_module/n33 [128]), 
            .CO(\test_module/add_41/n256 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i128 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i128 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i129  (.I0(o_pllBr0_reg[129]), .I1(1'b0), 
            .CI(\test_module/add_41/n256 ), .O(\test_module/n33 [129]), 
            .CO(\test_module/add_41/n258 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i129 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i129 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i130  (.I0(o_pllBr0_reg[130]), .I1(1'b0), 
            .CI(\test_module/add_41/n258 ), .O(\test_module/n33 [130]), 
            .CO(\test_module/add_41/n260 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i130 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i130 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i131  (.I0(o_pllBr0_reg[131]), .I1(1'b0), 
            .CI(\test_module/add_41/n260 ), .O(\test_module/n33 [131]), 
            .CO(\test_module/add_41/n262 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i131 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i131 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i132  (.I0(o_pllBr0_reg[132]), .I1(1'b0), 
            .CI(\test_module/add_41/n262 ), .O(\test_module/n33 [132]), 
            .CO(\test_module/add_41/n264 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i132 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i132 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i133  (.I0(o_pllBr0_reg[133]), .I1(1'b0), 
            .CI(\test_module/add_41/n264 ), .O(\test_module/n33 [133]), 
            .CO(\test_module/add_41/n266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i133 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i133 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i134  (.I0(o_pllBr0_reg[134]), .I1(1'b0), 
            .CI(\test_module/add_41/n266 ), .O(\test_module/n33 [134]), 
            .CO(\test_module/add_41/n268 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i134 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i134 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i135  (.I0(o_pllBr0_reg[135]), .I1(1'b0), 
            .CI(\test_module/add_41/n268 ), .O(\test_module/n33 [135]), 
            .CO(\test_module/add_41/n270 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i135 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i135 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i136  (.I0(o_pllBr0_reg[136]), .I1(1'b0), 
            .CI(\test_module/add_41/n270 ), .O(\test_module/n33 [136]), 
            .CO(\test_module/add_41/n272 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i136 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i136 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i137  (.I0(o_pllBr0_reg[137]), .I1(1'b0), 
            .CI(\test_module/add_41/n272 ), .O(\test_module/n33 [137]), 
            .CO(\test_module/add_41/n274 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i137 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i137 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i138  (.I0(o_pllBr0_reg[138]), .I1(1'b0), 
            .CI(\test_module/add_41/n274 ), .O(\test_module/n33 [138]), 
            .CO(\test_module/add_41/n276 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i138 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i138 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i139  (.I0(o_pllBr0_reg[139]), .I1(1'b0), 
            .CI(\test_module/add_41/n276 ), .O(\test_module/n33 [139]), 
            .CO(\test_module/add_41/n278 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i139 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i139 .I1_POLARITY = 1'b1;
    EFX_ADD \debug_inst/vio0/vio_core_inst/add_33/i2  (.I0(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I1(\debug_inst/vio0/vio_core_inst/opcode [1]), .CI(1'b0), .O(\debug_inst/vio0/vio_core_inst/incremented_address [1]), 
            .CO(\debug_inst/vio0/vio_core_inst/add_33/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1402)
    defparam \debug_inst/vio0/vio_core_inst/add_33/i2 .I0_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/add_33/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i66  (.I0(o_pllBr0_reg[66]), .I1(1'b0), 
            .CI(\test_module/add_41/n130 ), .O(\test_module/n33 [66]), .CO(\test_module/add_41/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i66 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i66 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i65  (.I0(o_pllBr0_reg[65]), .I1(1'b0), 
            .CI(\test_module/add_41/n128 ), .O(\test_module/n33 [65]), .CO(\test_module/add_41/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i65 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i65 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i89  (.I0(o_pllBr0_reg[89]), .I1(1'b0), 
            .CI(\test_module/add_41/n176 ), .O(\test_module/n33 [89]), .CO(\test_module/add_41/n178 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i89 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i89 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i92  (.I0(o_pllBr0_reg[92]), .I1(1'b0), 
            .CI(\test_module/add_41/n182 ), .O(\test_module/n33 [92]), .CO(\test_module/add_41/n184 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i92 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i92 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i140  (.I0(o_pllBr0_reg[140]), .I1(1'b0), 
            .CI(\test_module/add_41/n278 ), .O(\test_module/n33 [140]), 
            .CO(\test_module/add_41/n280 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i140 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i140 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i141  (.I0(o_pllBr0_reg[141]), .I1(1'b0), 
            .CI(\test_module/add_41/n280 ), .O(\test_module/n33 [141]), 
            .CO(\test_module/add_41/n282 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i141 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i141 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i142  (.I0(o_pllBr0_reg[142]), .I1(1'b0), 
            .CI(\test_module/add_41/n282 ), .O(\test_module/n33 [142]), 
            .CO(\test_module/add_41/n284 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i142 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i142 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i88  (.I0(o_pllBr0_reg[88]), .I1(1'b0), 
            .CI(\test_module/add_41/n174 ), .O(\test_module/n33 [88]), .CO(\test_module/add_41/n176 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i88 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i88 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i64  (.I0(o_pllBr0_reg[64]), .I1(1'b0), 
            .CI(\test_module/add_41/n126 ), .O(\test_module/n33 [64]), .CO(\test_module/add_41/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i64 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i64 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i63  (.I0(o_pllBr0_reg[63]), .I1(1'b0), 
            .CI(\test_module/add_41/n124 ), .O(\test_module/n33 [63]), .CO(\test_module/add_41/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i63 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i63 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i62  (.I0(o_pllBr0_reg[62]), .I1(1'b0), 
            .CI(\test_module/add_41/n122 ), .O(\test_module/n33 [62]), .CO(\test_module/add_41/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i62 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i62 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i61  (.I0(o_pllBr0_reg[61]), .I1(1'b0), 
            .CI(\test_module/add_41/n120 ), .O(\test_module/n33 [61]), .CO(\test_module/add_41/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i61 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i61 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i60  (.I0(o_pllBr0_reg[60]), .I1(1'b0), 
            .CI(\test_module/add_41/n118 ), .O(\test_module/n33 [60]), .CO(\test_module/add_41/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i60 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i60 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i59  (.I0(o_pllBr0_reg[59]), .I1(1'b0), 
            .CI(\test_module/add_41/n116 ), .O(\test_module/n33 [59]), .CO(\test_module/add_41/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i59 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i59 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i58  (.I0(o_pllBr0_reg[58]), .I1(1'b0), 
            .CI(\test_module/add_41/n114 ), .O(\test_module/n33 [58]), .CO(\test_module/add_41/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i58 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i58 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i57  (.I0(o_pllBr0_reg[57]), .I1(1'b0), 
            .CI(\test_module/add_41/n112 ), .O(\test_module/n33 [57]), .CO(\test_module/add_41/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i57 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i57 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i56  (.I0(o_pllBr0_reg[56]), .I1(1'b0), 
            .CI(\test_module/add_41/n110 ), .O(\test_module/n33 [56]), .CO(\test_module/add_41/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i56 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i56 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i55  (.I0(o_pllBr0_reg[55]), .I1(1'b0), 
            .CI(\test_module/add_41/n108 ), .O(\test_module/n33 [55]), .CO(\test_module/add_41/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i55 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i55 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i54  (.I0(o_pllBr0_reg[54]), .I1(1'b0), 
            .CI(\test_module/add_41/n106 ), .O(\test_module/n33 [54]), .CO(\test_module/add_41/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i54 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i54 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i53  (.I0(o_pllBr0_reg[53]), .I1(1'b0), 
            .CI(\test_module/add_41/n104 ), .O(\test_module/n33 [53]), .CO(\test_module/add_41/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i53 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i53 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i52  (.I0(o_pllBr0_reg[52]), .I1(1'b0), 
            .CI(\test_module/add_41/n102 ), .O(\test_module/n33 [52]), .CO(\test_module/add_41/n104 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i52 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i52 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i51  (.I0(o_pllBr0_reg[51]), .I1(1'b0), 
            .CI(\test_module/add_41/n100 ), .O(\test_module/n33 [51]), .CO(\test_module/add_41/n102 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i51 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i51 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i143  (.I0(o_pllBr0_reg[143]), .I1(1'b0), 
            .CI(\test_module/add_41/n284 ), .O(\test_module/n33 [143]), 
            .CO(\test_module/add_41/n286 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i143 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i143 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i144  (.I0(o_pllBr0_reg[144]), .I1(1'b0), 
            .CI(\test_module/add_41/n286 ), .O(\test_module/n33 [144]), 
            .CO(\test_module/add_41/n288 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i144 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i144 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i145  (.I0(o_pllBr0_reg[145]), .I1(1'b0), 
            .CI(\test_module/add_41/n288 ), .O(\test_module/n33 [145]), 
            .CO(\test_module/add_41/n290 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i145 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i145 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i146  (.I0(o_pllBr0_reg[146]), .I1(1'b0), 
            .CI(\test_module/add_41/n290 ), .O(\test_module/n33 [146]), 
            .CO(\test_module/add_41/n292 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i146 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i146 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i147  (.I0(o_pllBr0_reg[147]), .I1(1'b0), 
            .CI(\test_module/add_41/n292 ), .O(\test_module/n33 [147]), 
            .CO(\test_module/add_41/n294 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i147 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i147 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i148  (.I0(o_pllBr0_reg[148]), .I1(1'b0), 
            .CI(\test_module/add_41/n294 ), .O(\test_module/n33 [148]), 
            .CO(\test_module/add_41/n296 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i148 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i148 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i149  (.I0(o_pllBr0_reg[149]), .I1(1'b0), 
            .CI(\test_module/add_41/n296 ), .O(\test_module/n33 [149]), 
            .CO(\test_module/add_41/n298 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i149 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i149 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i150  (.I0(o_pllBr0_reg[150]), .I1(1'b0), 
            .CI(\test_module/add_41/n298 ), .O(\test_module/n33 [150]), 
            .CO(\test_module/add_41/n300 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i150 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i150 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i151  (.I0(o_pllBr0_reg[151]), .I1(1'b0), 
            .CI(\test_module/add_41/n300 ), .O(\test_module/n33 [151]), 
            .CO(\test_module/add_41/n302 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i151 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i151 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i152  (.I0(o_pllBr0_reg[152]), .I1(1'b0), 
            .CI(\test_module/add_41/n302 ), .O(\test_module/n33 [152]), 
            .CO(\test_module/add_41/n304 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i152 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i152 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i153  (.I0(o_pllBr0_reg[153]), .I1(1'b0), 
            .CI(\test_module/add_41/n304 ), .O(\test_module/n33 [153]), 
            .CO(\test_module/add_41/n306 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i153 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i153 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i154  (.I0(o_pllBr0_reg[154]), .I1(1'b0), 
            .CI(\test_module/add_41/n306 ), .O(\test_module/n33 [154]), 
            .CO(\test_module/add_41/n308 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i154 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i154 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i155  (.I0(o_pllBr0_reg[155]), .I1(1'b0), 
            .CI(\test_module/add_41/n308 ), .O(\test_module/n33 [155]), 
            .CO(\test_module/add_41/n310 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i155 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i155 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i156  (.I0(o_pllBr0_reg[156]), .I1(1'b0), 
            .CI(\test_module/add_41/n310 ), .O(\test_module/n33 [156]), 
            .CO(\test_module/add_41/n312 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i156 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i156 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i157  (.I0(o_pllBr0_reg[157]), .I1(1'b0), 
            .CI(\test_module/add_41/n312 ), .O(\test_module/n33 [157]), 
            .CO(\test_module/add_41/n314 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i157 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i157 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i158  (.I0(o_pllBr0_reg[158]), .I1(1'b0), 
            .CI(\test_module/add_41/n314 ), .O(\test_module/n33 [158]), 
            .CO(\test_module/add_41/n316 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i158 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i158 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i159  (.I0(o_pllBr0_reg[159]), .I1(1'b0), 
            .CI(\test_module/add_41/n316 ), .O(\test_module/n33 [159]), 
            .CO(\test_module/add_41/n318 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i159 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i159 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i160  (.I0(o_pllBr0_reg[160]), .I1(1'b0), 
            .CI(\test_module/add_41/n318 ), .O(\test_module/n33 [160]), 
            .CO(\test_module/add_41/n320 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i160 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i160 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i161  (.I0(o_pllBr0_reg[161]), .I1(1'b0), 
            .CI(\test_module/add_41/n320 ), .O(\test_module/n33 [161]), 
            .CO(\test_module/add_41/n322 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i161 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i161 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i162  (.I0(o_pllBr0_reg[162]), .I1(1'b0), 
            .CI(\test_module/add_41/n322 ), .O(\test_module/n33 [162]), 
            .CO(\test_module/add_41/n324 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i162 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i162 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i163  (.I0(o_pllBr0_reg[163]), .I1(1'b0), 
            .CI(\test_module/add_41/n324 ), .O(\test_module/n33 [163]), 
            .CO(\test_module/add_41/n326 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i163 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i163 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i164  (.I0(o_pllBr0_reg[164]), .I1(1'b0), 
            .CI(\test_module/add_41/n326 ), .O(\test_module/n33 [164]), 
            .CO(\test_module/add_41/n328 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i164 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i164 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i165  (.I0(o_pllBr0_reg[165]), .I1(1'b0), 
            .CI(\test_module/add_41/n328 ), .O(\test_module/n33 [165]), 
            .CO(\test_module/add_41/n330 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i165 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i165 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i166  (.I0(o_pllBr0_reg[166]), .I1(1'b0), 
            .CI(\test_module/add_41/n330 ), .O(\test_module/n33 [166]), 
            .CO(\test_module/add_41/n332 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i166 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i166 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i167  (.I0(o_pllBr0_reg[167]), .I1(1'b0), 
            .CI(\test_module/add_41/n332 ), .O(\test_module/n33 [167]), 
            .CO(\test_module/add_41/n334 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i167 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i167 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i168  (.I0(o_pllBr0_reg[168]), .I1(1'b0), 
            .CI(\test_module/add_41/n334 ), .O(\test_module/n33 [168]), 
            .CO(\test_module/add_41/n336 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i168 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i168 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i169  (.I0(o_pllBr0_reg[169]), .I1(1'b0), 
            .CI(\test_module/add_41/n336 ), .O(\test_module/n33 [169]), 
            .CO(\test_module/add_41/n338 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i169 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i169 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i170  (.I0(o_pllBr0_reg[170]), .I1(1'b0), 
            .CI(\test_module/add_41/n338 ), .O(\test_module/n33 [170]), 
            .CO(\test_module/add_41/n340 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i170 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i170 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i171  (.I0(o_pllBr0_reg[171]), .I1(1'b0), 
            .CI(\test_module/add_41/n340 ), .O(\test_module/n33 [171]), 
            .CO(\test_module/add_41/n342 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i171 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i171 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i172  (.I0(o_pllBr0_reg[172]), .I1(1'b0), 
            .CI(\test_module/add_41/n342 ), .O(\test_module/n33 [172]), 
            .CO(\test_module/add_41/n344 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i172 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i172 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i173  (.I0(o_pllBr0_reg[173]), .I1(1'b0), 
            .CI(\test_module/add_41/n344 ), .O(\test_module/n33 [173]), 
            .CO(\test_module/add_41/n346 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i173 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i173 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i174  (.I0(o_pllBr0_reg[174]), .I1(1'b0), 
            .CI(\test_module/add_41/n346 ), .O(\test_module/n33 [174]), 
            .CO(\test_module/add_41/n348 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i174 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i174 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i175  (.I0(o_pllBr0_reg[175]), .I1(1'b0), 
            .CI(\test_module/add_41/n348 ), .O(\test_module/n33 [175]), 
            .CO(\test_module/add_41/n350 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i175 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i175 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i176  (.I0(o_pllBr0_reg[176]), .I1(1'b0), 
            .CI(\test_module/add_41/n350 ), .O(\test_module/n33 [176]), 
            .CO(\test_module/add_41/n352 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i176 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i176 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i177  (.I0(o_pllBr0_reg[177]), .I1(1'b0), 
            .CI(\test_module/add_41/n352 ), .O(\test_module/n33 [177]), 
            .CO(\test_module/add_41/n354 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i177 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i177 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i178  (.I0(o_pllBr0_reg[178]), .I1(1'b0), 
            .CI(\test_module/add_41/n354 ), .O(\test_module/n33 [178]), 
            .CO(\test_module/add_41/n356 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i178 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i178 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i179  (.I0(o_pllBr0_reg[179]), .I1(1'b0), 
            .CI(\test_module/add_41/n356 ), .O(\test_module/n33 [179]), 
            .CO(\test_module/add_41/n358 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i179 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i179 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i180  (.I0(o_pllBr0_reg[180]), .I1(1'b0), 
            .CI(\test_module/add_41/n358 ), .O(\test_module/n33 [180]), 
            .CO(\test_module/add_41/n360 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i180 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i180 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i181  (.I0(o_pllBr0_reg[181]), .I1(1'b0), 
            .CI(\test_module/add_41/n360 ), .O(\test_module/n33 [181]), 
            .CO(\test_module/add_41/n362 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i181 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i181 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i182  (.I0(o_pllBr0_reg[182]), .I1(1'b0), 
            .CI(\test_module/add_41/n362 ), .O(\test_module/n33 [182]), 
            .CO(\test_module/add_41/n364 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i182 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i182 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i183  (.I0(o_pllBr0_reg[183]), .I1(1'b0), 
            .CI(\test_module/add_41/n364 ), .O(\test_module/n33 [183]), 
            .CO(\test_module/add_41/n366 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i183 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i183 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i184  (.I0(o_pllBr0_reg[184]), .I1(1'b0), 
            .CI(\test_module/add_41/n366 ), .O(\test_module/n33 [184]), 
            .CO(\test_module/add_41/n368 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i184 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i184 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i185  (.I0(o_pllBr0_reg[185]), .I1(1'b0), 
            .CI(\test_module/add_41/n368 ), .O(\test_module/n33 [185]), 
            .CO(\test_module/add_41/n370 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i185 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i185 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i186  (.I0(o_pllBr0_reg[186]), .I1(1'b0), 
            .CI(\test_module/add_41/n370 ), .O(\test_module/n33 [186]), 
            .CO(\test_module/add_41/n372 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i186 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i186 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i187  (.I0(o_pllBr0_reg[187]), .I1(1'b0), 
            .CI(\test_module/add_41/n372 ), .O(\test_module/n33 [187]), 
            .CO(\test_module/add_41/n374 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i187 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i187 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i188  (.I0(o_pllBr0_reg[188]), .I1(1'b0), 
            .CI(\test_module/add_41/n374 ), .O(\test_module/n33 [188]), 
            .CO(\test_module/add_41/n376 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i188 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i188 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i189  (.I0(o_pllBr0_reg[189]), .I1(1'b0), 
            .CI(\test_module/add_41/n376 ), .O(\test_module/n33 [189]), 
            .CO(\test_module/add_41/n378 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i189 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i189 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i190  (.I0(o_pllBr0_reg[190]), .I1(1'b0), 
            .CI(\test_module/add_41/n378 ), .O(\test_module/n33 [190]), 
            .CO(\test_module/add_41/n380 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i190 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i190 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i191  (.I0(o_pllBr0_reg[191]), .I1(1'b0), 
            .CI(\test_module/add_41/n380 ), .O(\test_module/n33 [191]), 
            .CO(\test_module/add_41/n382 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i191 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i191 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i192  (.I0(o_pllBr0_reg[192]), .I1(1'b0), 
            .CI(\test_module/add_41/n382 ), .O(\test_module/n33 [192]), 
            .CO(\test_module/add_41/n384 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i192 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i192 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i193  (.I0(o_pllBr0_reg[193]), .I1(1'b0), 
            .CI(\test_module/add_41/n384 ), .O(\test_module/n33 [193]), 
            .CO(\test_module/add_41/n386 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i193 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i193 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i194  (.I0(o_pllBr0_reg[194]), .I1(1'b0), 
            .CI(\test_module/add_41/n386 ), .O(\test_module/n33 [194]), 
            .CO(\test_module/add_41/n388 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i194 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i194 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i195  (.I0(o_pllBr0_reg[195]), .I1(1'b0), 
            .CI(\test_module/add_41/n388 ), .O(\test_module/n33 [195]), 
            .CO(\test_module/add_41/n390 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i195 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i195 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i196  (.I0(o_pllBr0_reg[196]), .I1(1'b0), 
            .CI(\test_module/add_41/n390 ), .O(\test_module/n33 [196]), 
            .CO(\test_module/add_41/n392 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i196 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i196 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i197  (.I0(o_pllBr0_reg[197]), .I1(1'b0), 
            .CI(\test_module/add_41/n392 ), .O(\test_module/n33 [197]), 
            .CO(\test_module/add_41/n394 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i197 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i197 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i198  (.I0(o_pllBr0_reg[198]), .I1(1'b0), 
            .CI(\test_module/add_41/n394 ), .O(\test_module/n33 [198]), 
            .CO(\test_module/add_41/n396 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i198 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i198 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i199  (.I0(o_pllBr0_reg[199]), .I1(1'b0), 
            .CI(\test_module/add_41/n396 ), .O(\test_module/n33 [199]), 
            .CO(\test_module/add_41/n398 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i199 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i199 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i200  (.I0(o_pllBr0_reg[200]), .I1(1'b0), 
            .CI(\test_module/add_41/n398 ), .O(\test_module/n33 [200]), 
            .CO(\test_module/add_41/n400 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i200 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i200 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i201  (.I0(o_pllBr0_reg[201]), .I1(1'b0), 
            .CI(\test_module/add_41/n400 ), .O(\test_module/n33 [201]), 
            .CO(\test_module/add_41/n402 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i201 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i201 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i202  (.I0(o_pllBr0_reg[202]), .I1(1'b0), 
            .CI(\test_module/add_41/n402 ), .O(\test_module/n33 [202]), 
            .CO(\test_module/add_41/n404 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i202 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i202 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i203  (.I0(o_pllBr0_reg[203]), .I1(1'b0), 
            .CI(\test_module/add_41/n404 ), .O(\test_module/n33 [203]), 
            .CO(\test_module/add_41/n406 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i203 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i203 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i204  (.I0(o_pllBr0_reg[204]), .I1(1'b0), 
            .CI(\test_module/add_41/n406 ), .O(\test_module/n33 [204]), 
            .CO(\test_module/add_41/n408 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i204 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i204 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i205  (.I0(o_pllBr0_reg[205]), .I1(1'b0), 
            .CI(\test_module/add_41/n408 ), .O(\test_module/n33 [205]), 
            .CO(\test_module/add_41/n410 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i205 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i205 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i206  (.I0(o_pllBr0_reg[206]), .I1(1'b0), 
            .CI(\test_module/add_41/n410 ), .O(\test_module/n33 [206]), 
            .CO(\test_module/add_41/n412 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i206 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i206 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i207  (.I0(o_pllBr0_reg[207]), .I1(1'b0), 
            .CI(\test_module/add_41/n412 ), .O(\test_module/n33 [207]), 
            .CO(\test_module/add_41/n414 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i207 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i207 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i208  (.I0(o_pllBr0_reg[208]), .I1(1'b0), 
            .CI(\test_module/add_41/n414 ), .O(\test_module/n33 [208]), 
            .CO(\test_module/add_41/n416 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i208 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i208 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i209  (.I0(o_pllBr0_reg[209]), .I1(1'b0), 
            .CI(\test_module/add_41/n416 ), .O(\test_module/n33 [209]), 
            .CO(\test_module/add_41/n418 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i209 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i209 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i210  (.I0(o_pllBr0_reg[210]), .I1(1'b0), 
            .CI(\test_module/add_41/n418 ), .O(\test_module/n33 [210]), 
            .CO(\test_module/add_41/n420 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i210 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i210 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i211  (.I0(o_pllBr0_reg[211]), .I1(1'b0), 
            .CI(\test_module/add_41/n420 ), .O(\test_module/n33 [211]), 
            .CO(\test_module/add_41/n422 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i211 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i211 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i212  (.I0(o_pllBr0_reg[212]), .I1(1'b0), 
            .CI(\test_module/add_41/n422 ), .O(\test_module/n33 [212]), 
            .CO(\test_module/add_41/n424 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i212 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i212 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i213  (.I0(o_pllBr0_reg[213]), .I1(1'b0), 
            .CI(\test_module/add_41/n424 ), .O(\test_module/n33 [213]), 
            .CO(\test_module/add_41/n426 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i213 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i213 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i214  (.I0(o_pllBr0_reg[214]), .I1(1'b0), 
            .CI(\test_module/add_41/n426 ), .O(\test_module/n33 [214]), 
            .CO(\test_module/add_41/n428 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i214 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i214 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i215  (.I0(o_pllBr0_reg[215]), .I1(1'b0), 
            .CI(\test_module/add_41/n428 ), .O(\test_module/n33 [215]), 
            .CO(\test_module/add_41/n430 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i215 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i215 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i216  (.I0(o_pllBr0_reg[216]), .I1(1'b0), 
            .CI(\test_module/add_41/n430 ), .O(\test_module/n33 [216]), 
            .CO(\test_module/add_41/n432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i216 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i216 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i217  (.I0(o_pllBr0_reg[217]), .I1(1'b0), 
            .CI(\test_module/add_41/n432 ), .O(\test_module/n33 [217]), 
            .CO(\test_module/add_41/n434 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i217 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i217 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i218  (.I0(o_pllBr0_reg[218]), .I1(1'b0), 
            .CI(\test_module/add_41/n434 ), .O(\test_module/n33 [218]), 
            .CO(\test_module/add_41/n436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i218 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i218 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i219  (.I0(o_pllBr0_reg[219]), .I1(1'b0), 
            .CI(\test_module/add_41/n436 ), .O(\test_module/n33 [219]), 
            .CO(\test_module/add_41/n438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i219 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i219 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i220  (.I0(o_pllBr0_reg[220]), .I1(1'b0), 
            .CI(\test_module/add_41/n438 ), .O(\test_module/n33 [220]), 
            .CO(\test_module/add_41/n440 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i220 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i220 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i221  (.I0(o_pllBr0_reg[221]), .I1(1'b0), 
            .CI(\test_module/add_41/n440 ), .O(\test_module/n33 [221]), 
            .CO(\test_module/add_41/n442 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i221 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i221 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i222  (.I0(o_pllBr0_reg[222]), .I1(1'b0), 
            .CI(\test_module/add_41/n442 ), .O(\test_module/n33 [222]), 
            .CO(\test_module/add_41/n444 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i222 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i222 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i223  (.I0(o_pllBr0_reg[223]), .I1(1'b0), 
            .CI(\test_module/add_41/n444 ), .O(\test_module/n33 [223]), 
            .CO(\test_module/add_41/n446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i223 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i223 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i224  (.I0(o_pllBr0_reg[224]), .I1(1'b0), 
            .CI(\test_module/add_41/n446 ), .O(\test_module/n33 [224]), 
            .CO(\test_module/add_41/n448 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i224 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i224 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i225  (.I0(o_pllBr0_reg[225]), .I1(1'b0), 
            .CI(\test_module/add_41/n448 ), .O(\test_module/n33 [225]), 
            .CO(\test_module/add_41/n450 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i225 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i225 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i226  (.I0(o_pllBr0_reg[226]), .I1(1'b0), 
            .CI(\test_module/add_41/n450 ), .O(\test_module/n33 [226]), 
            .CO(\test_module/add_41/n452 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i226 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i226 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i227  (.I0(o_pllBr0_reg[227]), .I1(1'b0), 
            .CI(\test_module/add_41/n452 ), .O(\test_module/n33 [227]), 
            .CO(\test_module/add_41/n454 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i227 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i227 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i228  (.I0(o_pllBr0_reg[228]), .I1(1'b0), 
            .CI(\test_module/add_41/n454 ), .O(\test_module/n33 [228]), 
            .CO(\test_module/add_41/n456 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i228 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i228 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i229  (.I0(o_pllBr0_reg[229]), .I1(1'b0), 
            .CI(\test_module/add_41/n456 ), .O(\test_module/n33 [229]), 
            .CO(\test_module/add_41/n458 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i229 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i229 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i230  (.I0(o_pllBr0_reg[230]), .I1(1'b0), 
            .CI(\test_module/add_41/n458 ), .O(\test_module/n33 [230]), 
            .CO(\test_module/add_41/n460 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i230 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i230 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i231  (.I0(o_pllBr0_reg[231]), .I1(1'b0), 
            .CI(\test_module/add_41/n460 ), .O(\test_module/n33 [231]), 
            .CO(\test_module/add_41/n462 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i231 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i231 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i232  (.I0(o_pllBr0_reg[232]), .I1(1'b0), 
            .CI(\test_module/add_41/n462 ), .O(\test_module/n33 [232]), 
            .CO(\test_module/add_41/n464 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i232 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i232 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i233  (.I0(o_pllBr0_reg[233]), .I1(1'b0), 
            .CI(\test_module/add_41/n464 ), .O(\test_module/n33 [233]), 
            .CO(\test_module/add_41/n466 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i233 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i233 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i234  (.I0(o_pllBr0_reg[234]), .I1(1'b0), 
            .CI(\test_module/add_41/n466 ), .O(\test_module/n33 [234]), 
            .CO(\test_module/add_41/n468 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i234 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i234 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i235  (.I0(o_pllBr0_reg[235]), .I1(1'b0), 
            .CI(\test_module/add_41/n468 ), .O(\test_module/n33 [235]), 
            .CO(\test_module/add_41/n470 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i235 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i235 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i236  (.I0(o_pllBr0_reg[236]), .I1(1'b0), 
            .CI(\test_module/add_41/n470 ), .O(\test_module/n33 [236]), 
            .CO(\test_module/add_41/n472 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i236 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i236 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i237  (.I0(o_pllBr0_reg[237]), .I1(1'b0), 
            .CI(\test_module/add_41/n472 ), .O(\test_module/n33 [237]), 
            .CO(\test_module/add_41/n474 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i237 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i237 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i238  (.I0(o_pllBr0_reg[238]), .I1(1'b0), 
            .CI(\test_module/add_41/n474 ), .O(\test_module/n33 [238]), 
            .CO(\test_module/add_41/n476 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i238 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i238 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i239  (.I0(o_pllBr0_reg[239]), .I1(1'b0), 
            .CI(\test_module/add_41/n476 ), .O(\test_module/n33 [239]), 
            .CO(\test_module/add_41/n478 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i239 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i239 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i240  (.I0(o_pllBr0_reg[240]), .I1(1'b0), 
            .CI(\test_module/add_41/n478 ), .O(\test_module/n33 [240]), 
            .CO(\test_module/add_41/n480 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i240 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i240 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i241  (.I0(o_pllBr0_reg[241]), .I1(1'b0), 
            .CI(\test_module/add_41/n480 ), .O(\test_module/n33 [241]), 
            .CO(\test_module/add_41/n482 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i241 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i241 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i242  (.I0(o_pllBr0_reg[242]), .I1(1'b0), 
            .CI(\test_module/add_41/n482 ), .O(\test_module/n33 [242]), 
            .CO(\test_module/add_41/n484 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i242 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i242 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i243  (.I0(o_pllBr0_reg[243]), .I1(1'b0), 
            .CI(\test_module/add_41/n484 ), .O(\test_module/n33 [243]), 
            .CO(\test_module/add_41/n486 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i243 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i243 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i244  (.I0(o_pllBr0_reg[244]), .I1(1'b0), 
            .CI(\test_module/add_41/n486 ), .O(\test_module/n33 [244]), 
            .CO(\test_module/add_41/n488 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i244 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i244 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i245  (.I0(o_pllBr0_reg[245]), .I1(1'b0), 
            .CI(\test_module/add_41/n488 ), .O(\test_module/n33 [245]), 
            .CO(\test_module/add_41/n490 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i245 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i245 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i246  (.I0(o_pllBr0_reg[246]), .I1(1'b0), 
            .CI(\test_module/add_41/n490 ), .O(\test_module/n33 [246]), 
            .CO(\test_module/add_41/n492 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i246 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i246 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i247  (.I0(o_pllBr0_reg[247]), .I1(1'b0), 
            .CI(\test_module/add_41/n492 ), .O(\test_module/n33 [247]), 
            .CO(\test_module/add_41/n494 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i247 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i247 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i248  (.I0(o_pllBr0_reg[248]), .I1(1'b0), 
            .CI(\test_module/add_41/n494 ), .O(\test_module/n33 [248]), 
            .CO(\test_module/add_41/n496 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i248 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i248 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i249  (.I0(o_pllBr0_reg[249]), .I1(1'b0), 
            .CI(\test_module/add_41/n496 ), .O(\test_module/n33 [249]), 
            .CO(\test_module/add_41/n498 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i249 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i249 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i250  (.I0(o_pllBr0_reg[250]), .I1(1'b0), 
            .CI(\test_module/add_41/n498 ), .O(\test_module/n33 [250]), 
            .CO(\test_module/add_41/n500 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i250 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i250 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i251  (.I0(o_pllBr0_reg[251]), .I1(1'b0), 
            .CI(\test_module/add_41/n500 ), .O(\test_module/n33 [251]), 
            .CO(\test_module/add_41/n502 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i251 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i251 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i252  (.I0(o_pllBr0_reg[252]), .I1(1'b0), 
            .CI(\test_module/add_41/n502 ), .O(\test_module/n33 [252]), 
            .CO(\test_module/add_41/n504 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i252 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i252 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i253  (.I0(o_pllBr0_reg[253]), .I1(1'b0), 
            .CI(\test_module/add_41/n504 ), .O(\test_module/n33 [253]), 
            .CO(\test_module/add_41/n506 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i253 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i253 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i254  (.I0(o_pllBr0_reg[254]), .I1(1'b0), 
            .CI(\test_module/add_41/n506 ), .O(\test_module/n33 [254]), 
            .CO(\test_module/add_41/n508 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i254 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i254 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i255  (.I0(o_pllBr0_reg[255]), .I1(1'b0), 
            .CI(\test_module/add_41/n508 ), .O(\test_module/n33 [255])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i255 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i255 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_44/i2  (.I0(\test_module/delay_2 [2]), .I1(1'b0), 
            .CI(\test_module/add_44/n2 ), .O(\test_module/n1132 [2]), .CO(\test_module/add_44/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(34)
    defparam \test_module/add_44/i2 .I0_POLARITY = 1'b1;
    defparam \test_module/add_44/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_44/i3  (.I0(\test_module/delay_2 [3]), .I1(1'b0), 
            .CI(\test_module/add_44/n4 ), .O(\test_module/n1132 [3]), .CO(\test_module/add_44/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(34)
    defparam \test_module/add_44/i3 .I0_POLARITY = 1'b1;
    defparam \test_module/add_44/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_44/i4  (.I0(\test_module/delay_2 [4]), .I1(1'b0), 
            .CI(\test_module/add_44/n6 ), .O(\test_module/n1132 [4]), .CO(\test_module/add_44/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(34)
    defparam \test_module/add_44/i4 .I0_POLARITY = 1'b1;
    defparam \test_module/add_44/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_44/i5  (.I0(\test_module/delay_2 [5]), .I1(1'b0), 
            .CI(\test_module/add_44/n8 ), .O(\test_module/n1132 [5]), .CO(\test_module/add_44/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(34)
    defparam \test_module/add_44/i5 .I0_POLARITY = 1'b1;
    defparam \test_module/add_44/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_44/i6  (.I0(\test_module/delay_2 [6]), .I1(1'b0), 
            .CI(\test_module/add_44/n10 ), .O(\test_module/n1132 [6]), .CO(\test_module/add_44/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(34)
    defparam \test_module/add_44/i6 .I0_POLARITY = 1'b1;
    defparam \test_module/add_44/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_44/i7  (.I0(\test_module/delay_2 [7]), .I1(1'b0), 
            .CI(\test_module/add_44/n12 ), .O(\test_module/n1132 [7]), .CO(\test_module/add_44/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(34)
    defparam \test_module/add_44/i7 .I0_POLARITY = 1'b1;
    defparam \test_module/add_44/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_44/i8  (.I0(\test_module/delay_2 [8]), .I1(1'b0), 
            .CI(\test_module/add_44/n14 ), .O(\test_module/n1132 [8]), .CO(\test_module/add_44/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(34)
    defparam \test_module/add_44/i8 .I0_POLARITY = 1'b1;
    defparam \test_module/add_44/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_44/i9  (.I0(\test_module/delay_2 [9]), .I1(1'b0), 
            .CI(\test_module/add_44/n16 ), .O(\test_module/n1132 [9]), .CO(\test_module/add_44/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(34)
    defparam \test_module/add_44/i9 .I0_POLARITY = 1'b1;
    defparam \test_module/add_44/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_44/i10  (.I0(\test_module/delay_2 [10]), .I1(1'b0), 
            .CI(\test_module/add_44/n18 ), .O(\test_module/n1132 [10]), 
            .CO(\test_module/add_44/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(34)
    defparam \test_module/add_44/i10 .I0_POLARITY = 1'b1;
    defparam \test_module/add_44/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_44/i11  (.I0(\test_module/delay_2 [11]), .I1(1'b0), 
            .CI(\test_module/add_44/n20 ), .O(\test_module/n1132 [11]), 
            .CO(\test_module/add_44/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(34)
    defparam \test_module/add_44/i11 .I0_POLARITY = 1'b1;
    defparam \test_module/add_44/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_44/i12  (.I0(\test_module/delay_2 [12]), .I1(1'b0), 
            .CI(\test_module/add_44/n22 ), .O(\test_module/n1132 [12]), 
            .CO(\test_module/add_44/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(34)
    defparam \test_module/add_44/i12 .I0_POLARITY = 1'b1;
    defparam \test_module/add_44/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_44/i13  (.I0(\test_module/delay_2 [13]), .I1(1'b0), 
            .CI(\test_module/add_44/n24 ), .O(\test_module/n1132 [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(34)
    defparam \test_module/add_44/i13 .I0_POLARITY = 1'b1;
    defparam \test_module/add_44/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i2  (.I0(o_pllBr1_reg[2]), .I1(1'b0), .CI(\test_module/add_46/n2 ), 
            .O(\test_module/n1156 [2]), .CO(\test_module/add_46/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i2 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i3  (.I0(o_pllBr1_reg[3]), .I1(1'b0), .CI(\test_module/add_46/n4 ), 
            .O(\test_module/n1156 [3]), .CO(\test_module/add_46/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i3 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i4  (.I0(o_pllBr1_reg[4]), .I1(1'b0), .CI(\test_module/add_46/n6 ), 
            .O(\test_module/n1156 [4]), .CO(\test_module/add_46/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i4 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i5  (.I0(o_pllBr1_reg[5]), .I1(1'b0), .CI(\test_module/add_46/n8 ), 
            .O(\test_module/n1156 [5]), .CO(\test_module/add_46/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i5 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i6  (.I0(o_pllBr1_reg[6]), .I1(1'b0), .CI(\test_module/add_46/n10 ), 
            .O(\test_module/n1156 [6]), .CO(\test_module/add_46/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i6 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i7  (.I0(o_pllBr1_reg[7]), .I1(1'b0), .CI(\test_module/add_46/n12 ), 
            .O(\test_module/n1156 [7]), .CO(\test_module/add_46/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i7 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i8  (.I0(o_pllBr1_reg[8]), .I1(1'b0), .CI(\test_module/add_46/n14 ), 
            .O(\test_module/n1156 [8]), .CO(\test_module/add_46/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i8 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i9  (.I0(o_pllBr1_reg[9]), .I1(1'b0), .CI(\test_module/add_46/n16 ), 
            .O(\test_module/n1156 [9]), .CO(\test_module/add_46/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i9 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i10  (.I0(o_pllBr1_reg[10]), .I1(1'b0), 
            .CI(\test_module/add_46/n18 ), .O(\test_module/n1156 [10]), 
            .CO(\test_module/add_46/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i10 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i11  (.I0(o_pllBr1_reg[11]), .I1(1'b0), 
            .CI(\test_module/add_46/n20 ), .O(\test_module/n1156 [11]), 
            .CO(\test_module/add_46/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i11 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i12  (.I0(o_pllBr1_reg[12]), .I1(1'b0), 
            .CI(\test_module/add_46/n22 ), .O(\test_module/n1156 [12]), 
            .CO(\test_module/add_46/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i12 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i13  (.I0(o_pllBr1_reg[13]), .I1(1'b0), 
            .CI(\test_module/add_46/n24 ), .O(\test_module/n1156 [13]), 
            .CO(\test_module/add_46/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i13 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i14  (.I0(o_pllBr1_reg[14]), .I1(1'b0), 
            .CI(\test_module/add_46/n26 ), .O(\test_module/n1156 [14]), 
            .CO(\test_module/add_46/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i14 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i15  (.I0(o_pllBr1_reg[15]), .I1(1'b0), 
            .CI(\test_module/add_46/n28 ), .O(\test_module/n1156 [15]), 
            .CO(\test_module/add_46/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i15 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i16  (.I0(o_pllBr1_reg[16]), .I1(1'b0), 
            .CI(\test_module/add_46/n30 ), .O(\test_module/n1156 [16]), 
            .CO(\test_module/add_46/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i16 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i17  (.I0(o_pllBr1_reg[17]), .I1(1'b0), 
            .CI(\test_module/add_46/n32 ), .O(\test_module/n1156 [17]), 
            .CO(\test_module/add_46/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i17 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i18  (.I0(o_pllBr1_reg[18]), .I1(1'b0), 
            .CI(\test_module/add_46/n34 ), .O(\test_module/n1156 [18]), 
            .CO(\test_module/add_46/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i18 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i19  (.I0(o_pllBr1_reg[19]), .I1(1'b0), 
            .CI(\test_module/add_46/n36 ), .O(\test_module/n1156 [19]), 
            .CO(\test_module/add_46/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i19 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i20  (.I0(o_pllBr1_reg[20]), .I1(1'b0), 
            .CI(\test_module/add_46/n38 ), .O(\test_module/n1156 [20]), 
            .CO(\test_module/add_46/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i20 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i21  (.I0(o_pllBr1_reg[21]), .I1(1'b0), 
            .CI(\test_module/add_46/n40 ), .O(\test_module/n1156 [21]), 
            .CO(\test_module/add_46/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i21 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i22  (.I0(o_pllBr1_reg[22]), .I1(1'b0), 
            .CI(\test_module/add_46/n42 ), .O(\test_module/n1156 [22]), 
            .CO(\test_module/add_46/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i22 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i23  (.I0(o_pllBr1_reg[23]), .I1(1'b0), 
            .CI(\test_module/add_46/n44 ), .O(\test_module/n1156 [23]), 
            .CO(\test_module/add_46/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i23 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i24  (.I0(o_pllBr1_reg[24]), .I1(1'b0), 
            .CI(\test_module/add_46/n46 ), .O(\test_module/n1156 [24]), 
            .CO(\test_module/add_46/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i24 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i25  (.I0(o_pllBr1_reg[25]), .I1(1'b0), 
            .CI(\test_module/add_46/n48 ), .O(\test_module/n1156 [25]), 
            .CO(\test_module/add_46/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i25 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i26  (.I0(o_pllBr1_reg[26]), .I1(1'b0), 
            .CI(\test_module/add_46/n50 ), .O(\test_module/n1156 [26]), 
            .CO(\test_module/add_46/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i26 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i27  (.I0(o_pllBr1_reg[27]), .I1(1'b0), 
            .CI(\test_module/add_46/n52 ), .O(\test_module/n1156 [27]), 
            .CO(\test_module/add_46/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i27 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i28  (.I0(o_pllBr1_reg[28]), .I1(1'b0), 
            .CI(\test_module/add_46/n54 ), .O(\test_module/n1156 [28]), 
            .CO(\test_module/add_46/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i28 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i29  (.I0(o_pllBr1_reg[29]), .I1(1'b0), 
            .CI(\test_module/add_46/n56 ), .O(\test_module/n1156 [29]), 
            .CO(\test_module/add_46/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i29 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i30  (.I0(o_pllBr1_reg[30]), .I1(1'b0), 
            .CI(\test_module/add_46/n58 ), .O(\test_module/n1156 [30]), 
            .CO(\test_module/add_46/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i30 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i31  (.I0(o_pllBr1_reg[31]), .I1(1'b0), 
            .CI(\test_module/add_46/n60 ), .O(\test_module/n1156 [31]), 
            .CO(\test_module/add_46/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i31 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i32  (.I0(o_pllBr1_reg[32]), .I1(1'b0), 
            .CI(\test_module/add_46/n62 ), .O(\test_module/n1156 [32]), 
            .CO(\test_module/add_46/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i32 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i33  (.I0(o_pllBr1_reg[33]), .I1(1'b0), 
            .CI(\test_module/add_46/n64 ), .O(\test_module/n1156 [33]), 
            .CO(\test_module/add_46/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i33 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i33 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i34  (.I0(o_pllBr1_reg[34]), .I1(1'b0), 
            .CI(\test_module/add_46/n66 ), .O(\test_module/n1156 [34]), 
            .CO(\test_module/add_46/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i34 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i34 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i35  (.I0(o_pllBr1_reg[35]), .I1(1'b0), 
            .CI(\test_module/add_46/n68 ), .O(\test_module/n1156 [35]), 
            .CO(\test_module/add_46/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i35 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i35 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i36  (.I0(o_pllBr1_reg[36]), .I1(1'b0), 
            .CI(\test_module/add_46/n70 ), .O(\test_module/n1156 [36]), 
            .CO(\test_module/add_46/n72 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i36 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i36 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i37  (.I0(o_pllBr1_reg[37]), .I1(1'b0), 
            .CI(\test_module/add_46/n72 ), .O(\test_module/n1156 [37]), 
            .CO(\test_module/add_46/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i37 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i37 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i38  (.I0(o_pllBr1_reg[38]), .I1(1'b0), 
            .CI(\test_module/add_46/n74 ), .O(\test_module/n1156 [38]), 
            .CO(\test_module/add_46/n76 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i38 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i38 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i39  (.I0(o_pllBr1_reg[39]), .I1(1'b0), 
            .CI(\test_module/add_46/n76 ), .O(\test_module/n1156 [39]), 
            .CO(\test_module/add_46/n78 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i39 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i39 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i40  (.I0(o_pllBr1_reg[40]), .I1(1'b0), 
            .CI(\test_module/add_46/n78 ), .O(\test_module/n1156 [40]), 
            .CO(\test_module/add_46/n80 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i40 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i40 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i41  (.I0(o_pllBr1_reg[41]), .I1(1'b0), 
            .CI(\test_module/add_46/n80 ), .O(\test_module/n1156 [41]), 
            .CO(\test_module/add_46/n82 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i41 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i41 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i42  (.I0(o_pllBr1_reg[42]), .I1(1'b0), 
            .CI(\test_module/add_46/n82 ), .O(\test_module/n1156 [42]), 
            .CO(\test_module/add_46/n84 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i42 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i42 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i43  (.I0(o_pllBr1_reg[43]), .I1(1'b0), 
            .CI(\test_module/add_46/n84 ), .O(\test_module/n1156 [43]), 
            .CO(\test_module/add_46/n86 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i43 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i43 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i44  (.I0(o_pllBr1_reg[44]), .I1(1'b0), 
            .CI(\test_module/add_46/n86 ), .O(\test_module/n1156 [44]), 
            .CO(\test_module/add_46/n88 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i44 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i44 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i45  (.I0(o_pllBr1_reg[45]), .I1(1'b0), 
            .CI(\test_module/add_46/n88 ), .O(\test_module/n1156 [45]), 
            .CO(\test_module/add_46/n90 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i45 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i45 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i46  (.I0(o_pllBr1_reg[46]), .I1(1'b0), 
            .CI(\test_module/add_46/n90 ), .O(\test_module/n1156 [46]), 
            .CO(\test_module/add_46/n92 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i46 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i46 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i47  (.I0(o_pllBr1_reg[47]), .I1(1'b0), 
            .CI(\test_module/add_46/n92 ), .O(\test_module/n1156 [47]), 
            .CO(\test_module/add_46/n94 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i47 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i47 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i48  (.I0(o_pllBr1_reg[48]), .I1(1'b0), 
            .CI(\test_module/add_46/n94 ), .O(\test_module/n1156 [48]), 
            .CO(\test_module/add_46/n96 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i48 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i48 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i49  (.I0(o_pllBr1_reg[49]), .I1(1'b0), 
            .CI(\test_module/add_46/n96 ), .O(\test_module/n1156 [49]), 
            .CO(\test_module/add_46/n98 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i49 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i49 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i50  (.I0(o_pllBr1_reg[50]), .I1(1'b0), 
            .CI(\test_module/add_46/n98 ), .O(\test_module/n1156 [50]), 
            .CO(\test_module/add_46/n100 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i50 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i50 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i51  (.I0(o_pllBr1_reg[51]), .I1(1'b0), 
            .CI(\test_module/add_46/n100 ), .O(\test_module/n1156 [51]), 
            .CO(\test_module/add_46/n102 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i51 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i51 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i52  (.I0(o_pllBr1_reg[52]), .I1(1'b0), 
            .CI(\test_module/add_46/n102 ), .O(\test_module/n1156 [52]), 
            .CO(\test_module/add_46/n104 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i52 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i52 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i53  (.I0(o_pllBr1_reg[53]), .I1(1'b0), 
            .CI(\test_module/add_46/n104 ), .O(\test_module/n1156 [53]), 
            .CO(\test_module/add_46/n106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i53 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i53 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i54  (.I0(o_pllBr1_reg[54]), .I1(1'b0), 
            .CI(\test_module/add_46/n106 ), .O(\test_module/n1156 [54]), 
            .CO(\test_module/add_46/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i54 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i54 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i55  (.I0(o_pllBr1_reg[55]), .I1(1'b0), 
            .CI(\test_module/add_46/n108 ), .O(\test_module/n1156 [55]), 
            .CO(\test_module/add_46/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i55 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i55 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i56  (.I0(o_pllBr1_reg[56]), .I1(1'b0), 
            .CI(\test_module/add_46/n110 ), .O(\test_module/n1156 [56]), 
            .CO(\test_module/add_46/n112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i56 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i56 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i57  (.I0(o_pllBr1_reg[57]), .I1(1'b0), 
            .CI(\test_module/add_46/n112 ), .O(\test_module/n1156 [57]), 
            .CO(\test_module/add_46/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i57 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i57 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i58  (.I0(o_pllBr1_reg[58]), .I1(1'b0), 
            .CI(\test_module/add_46/n114 ), .O(\test_module/n1156 [58]), 
            .CO(\test_module/add_46/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i58 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i58 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i59  (.I0(o_pllBr1_reg[59]), .I1(1'b0), 
            .CI(\test_module/add_46/n116 ), .O(\test_module/n1156 [59]), 
            .CO(\test_module/add_46/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i59 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i59 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i60  (.I0(o_pllBr1_reg[60]), .I1(1'b0), 
            .CI(\test_module/add_46/n118 ), .O(\test_module/n1156 [60]), 
            .CO(\test_module/add_46/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i60 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i60 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i61  (.I0(o_pllBr1_reg[61]), .I1(1'b0), 
            .CI(\test_module/add_46/n120 ), .O(\test_module/n1156 [61]), 
            .CO(\test_module/add_46/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i61 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i61 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i62  (.I0(o_pllBr1_reg[62]), .I1(1'b0), 
            .CI(\test_module/add_46/n122 ), .O(\test_module/n1156 [62]), 
            .CO(\test_module/add_46/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i62 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i62 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i63  (.I0(o_pllBr1_reg[63]), .I1(1'b0), 
            .CI(\test_module/add_46/n124 ), .O(\test_module/n1156 [63]), 
            .CO(\test_module/add_46/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i63 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i63 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i64  (.I0(o_pllBr1_reg[64]), .I1(1'b0), 
            .CI(\test_module/add_46/n126 ), .O(\test_module/n1156 [64]), 
            .CO(\test_module/add_46/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i64 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i64 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i65  (.I0(o_pllBr1_reg[65]), .I1(1'b0), 
            .CI(\test_module/add_46/n128 ), .O(\test_module/n1156 [65]), 
            .CO(\test_module/add_46/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i65 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i65 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i66  (.I0(o_pllBr1_reg[66]), .I1(1'b0), 
            .CI(\test_module/add_46/n130 ), .O(\test_module/n1156 [66]), 
            .CO(\test_module/add_46/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i66 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i66 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i67  (.I0(o_pllBr1_reg[67]), .I1(1'b0), 
            .CI(\test_module/add_46/n132 ), .O(\test_module/n1156 [67]), 
            .CO(\test_module/add_46/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i67 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i67 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i68  (.I0(o_pllBr1_reg[68]), .I1(1'b0), 
            .CI(\test_module/add_46/n134 ), .O(\test_module/n1156 [68]), 
            .CO(\test_module/add_46/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i68 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i68 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i69  (.I0(o_pllBr1_reg[69]), .I1(1'b0), 
            .CI(\test_module/add_46/n136 ), .O(\test_module/n1156 [69]), 
            .CO(\test_module/add_46/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i69 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i69 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i70  (.I0(o_pllBr1_reg[70]), .I1(1'b0), 
            .CI(\test_module/add_46/n138 ), .O(\test_module/n1156 [70]), 
            .CO(\test_module/add_46/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i70 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i70 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i71  (.I0(o_pllBr1_reg[71]), .I1(1'b0), 
            .CI(\test_module/add_46/n140 ), .O(\test_module/n1156 [71]), 
            .CO(\test_module/add_46/n142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i71 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i71 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i72  (.I0(o_pllBr1_reg[72]), .I1(1'b0), 
            .CI(\test_module/add_46/n142 ), .O(\test_module/n1156 [72]), 
            .CO(\test_module/add_46/n144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i72 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i72 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i73  (.I0(o_pllBr1_reg[73]), .I1(1'b0), 
            .CI(\test_module/add_46/n144 ), .O(\test_module/n1156 [73]), 
            .CO(\test_module/add_46/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i73 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i73 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i74  (.I0(o_pllBr1_reg[74]), .I1(1'b0), 
            .CI(\test_module/add_46/n146 ), .O(\test_module/n1156 [74]), 
            .CO(\test_module/add_46/n148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i74 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i74 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i75  (.I0(o_pllBr1_reg[75]), .I1(1'b0), 
            .CI(\test_module/add_46/n148 ), .O(\test_module/n1156 [75]), 
            .CO(\test_module/add_46/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i75 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i75 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i76  (.I0(o_pllBr1_reg[76]), .I1(1'b0), 
            .CI(\test_module/add_46/n150 ), .O(\test_module/n1156 [76]), 
            .CO(\test_module/add_46/n152 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i76 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i76 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i77  (.I0(o_pllBr1_reg[77]), .I1(1'b0), 
            .CI(\test_module/add_46/n152 ), .O(\test_module/n1156 [77]), 
            .CO(\test_module/add_46/n154 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i77 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i77 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i78  (.I0(o_pllBr1_reg[78]), .I1(1'b0), 
            .CI(\test_module/add_46/n154 ), .O(\test_module/n1156 [78]), 
            .CO(\test_module/add_46/n156 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i78 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i78 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i79  (.I0(o_pllBr1_reg[79]), .I1(1'b0), 
            .CI(\test_module/add_46/n156 ), .O(\test_module/n1156 [79]), 
            .CO(\test_module/add_46/n158 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i79 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i79 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i80  (.I0(o_pllBr1_reg[80]), .I1(1'b0), 
            .CI(\test_module/add_46/n158 ), .O(\test_module/n1156 [80]), 
            .CO(\test_module/add_46/n160 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i80 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i80 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i81  (.I0(o_pllBr1_reg[81]), .I1(1'b0), 
            .CI(\test_module/add_46/n160 ), .O(\test_module/n1156 [81]), 
            .CO(\test_module/add_46/n162 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i81 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i81 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i82  (.I0(o_pllBr1_reg[82]), .I1(1'b0), 
            .CI(\test_module/add_46/n162 ), .O(\test_module/n1156 [82]), 
            .CO(\test_module/add_46/n164 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i82 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i82 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i83  (.I0(o_pllBr1_reg[83]), .I1(1'b0), 
            .CI(\test_module/add_46/n164 ), .O(\test_module/n1156 [83]), 
            .CO(\test_module/add_46/n166 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i83 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i83 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i84  (.I0(o_pllBr1_reg[84]), .I1(1'b0), 
            .CI(\test_module/add_46/n166 ), .O(\test_module/n1156 [84]), 
            .CO(\test_module/add_46/n168 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i84 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i84 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i85  (.I0(o_pllBr1_reg[85]), .I1(1'b0), 
            .CI(\test_module/add_46/n168 ), .O(\test_module/n1156 [85]), 
            .CO(\test_module/add_46/n170 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i85 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i85 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i86  (.I0(o_pllBr1_reg[86]), .I1(1'b0), 
            .CI(\test_module/add_46/n170 ), .O(\test_module/n1156 [86]), 
            .CO(\test_module/add_46/n172 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i86 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i86 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i87  (.I0(o_pllBr1_reg[87]), .I1(1'b0), 
            .CI(\test_module/add_46/n172 ), .O(\test_module/n1156 [87]), 
            .CO(\test_module/add_46/n174 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i87 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i87 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i88  (.I0(o_pllBr1_reg[88]), .I1(1'b0), 
            .CI(\test_module/add_46/n174 ), .O(\test_module/n1156 [88]), 
            .CO(\test_module/add_46/n176 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i88 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i88 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i89  (.I0(o_pllBr1_reg[89]), .I1(1'b0), 
            .CI(\test_module/add_46/n176 ), .O(\test_module/n1156 [89]), 
            .CO(\test_module/add_46/n178 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i89 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i89 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i90  (.I0(o_pllBr1_reg[90]), .I1(1'b0), 
            .CI(\test_module/add_46/n178 ), .O(\test_module/n1156 [90]), 
            .CO(\test_module/add_46/n180 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i90 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i90 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i91  (.I0(o_pllBr1_reg[91]), .I1(1'b0), 
            .CI(\test_module/add_46/n180 ), .O(\test_module/n1156 [91]), 
            .CO(\test_module/add_46/n182 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i91 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i91 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i92  (.I0(o_pllBr1_reg[92]), .I1(1'b0), 
            .CI(\test_module/add_46/n182 ), .O(\test_module/n1156 [92]), 
            .CO(\test_module/add_46/n184 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i92 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i92 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i93  (.I0(o_pllBr1_reg[93]), .I1(1'b0), 
            .CI(\test_module/add_46/n184 ), .O(\test_module/n1156 [93]), 
            .CO(\test_module/add_46/n186 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i93 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i93 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i94  (.I0(o_pllBr1_reg[94]), .I1(1'b0), 
            .CI(\test_module/add_46/n186 ), .O(\test_module/n1156 [94]), 
            .CO(\test_module/add_46/n188 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i94 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i94 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i95  (.I0(o_pllBr1_reg[95]), .I1(1'b0), 
            .CI(\test_module/add_46/n188 ), .O(\test_module/n1156 [95]), 
            .CO(\test_module/add_46/n190 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i95 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i95 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i96  (.I0(o_pllBr1_reg[96]), .I1(1'b0), 
            .CI(\test_module/add_46/n190 ), .O(\test_module/n1156 [96]), 
            .CO(\test_module/add_46/n192 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i96 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i96 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i97  (.I0(o_pllBr1_reg[97]), .I1(1'b0), 
            .CI(\test_module/add_46/n192 ), .O(\test_module/n1156 [97]), 
            .CO(\test_module/add_46/n194 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i97 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i97 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i98  (.I0(o_pllBr1_reg[98]), .I1(1'b0), 
            .CI(\test_module/add_46/n194 ), .O(\test_module/n1156 [98]), 
            .CO(\test_module/add_46/n196 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i98 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i98 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i99  (.I0(o_pllBr1_reg[99]), .I1(1'b0), 
            .CI(\test_module/add_46/n196 ), .O(\test_module/n1156 [99]), 
            .CO(\test_module/add_46/n198 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i99 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i99 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i100  (.I0(o_pllBr1_reg[100]), .I1(1'b0), 
            .CI(\test_module/add_46/n198 ), .O(\test_module/n1156 [100]), 
            .CO(\test_module/add_46/n200 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i100 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i100 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i101  (.I0(o_pllBr1_reg[101]), .I1(1'b0), 
            .CI(\test_module/add_46/n200 ), .O(\test_module/n1156 [101]), 
            .CO(\test_module/add_46/n202 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i101 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i101 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i102  (.I0(o_pllBr1_reg[102]), .I1(1'b0), 
            .CI(\test_module/add_46/n202 ), .O(\test_module/n1156 [102]), 
            .CO(\test_module/add_46/n204 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i102 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i102 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i103  (.I0(o_pllBr1_reg[103]), .I1(1'b0), 
            .CI(\test_module/add_46/n204 ), .O(\test_module/n1156 [103]), 
            .CO(\test_module/add_46/n206 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i103 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i103 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i104  (.I0(o_pllBr1_reg[104]), .I1(1'b0), 
            .CI(\test_module/add_46/n206 ), .O(\test_module/n1156 [104]), 
            .CO(\test_module/add_46/n208 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i104 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i104 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i105  (.I0(o_pllBr1_reg[105]), .I1(1'b0), 
            .CI(\test_module/add_46/n208 ), .O(\test_module/n1156 [105]), 
            .CO(\test_module/add_46/n210 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i105 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i105 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i106  (.I0(o_pllBr1_reg[106]), .I1(1'b0), 
            .CI(\test_module/add_46/n210 ), .O(\test_module/n1156 [106]), 
            .CO(\test_module/add_46/n212 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i106 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i106 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i107  (.I0(o_pllBr1_reg[107]), .I1(1'b0), 
            .CI(\test_module/add_46/n212 ), .O(\test_module/n1156 [107]), 
            .CO(\test_module/add_46/n214 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i107 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i107 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i108  (.I0(o_pllBr1_reg[108]), .I1(1'b0), 
            .CI(\test_module/add_46/n214 ), .O(\test_module/n1156 [108]), 
            .CO(\test_module/add_46/n216 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i108 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i108 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i109  (.I0(o_pllBr1_reg[109]), .I1(1'b0), 
            .CI(\test_module/add_46/n216 ), .O(\test_module/n1156 [109]), 
            .CO(\test_module/add_46/n218 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i109 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i109 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i91  (.I0(o_pllBr0_reg[91]), .I1(1'b0), 
            .CI(\test_module/add_41/n180 ), .O(\test_module/n33 [91]), .CO(\test_module/add_41/n182 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i91 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i91 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i110  (.I0(o_pllBr1_reg[110]), .I1(1'b0), 
            .CI(\test_module/add_46/n218 ), .O(\test_module/n1156 [110]), 
            .CO(\test_module/add_46/n220 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i110 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i110 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i111  (.I0(o_pllBr1_reg[111]), .I1(1'b0), 
            .CI(\test_module/add_46/n220 ), .O(\test_module/n1156 [111]), 
            .CO(\test_module/add_46/n222 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i111 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i111 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i112  (.I0(o_pllBr1_reg[112]), .I1(1'b0), 
            .CI(\test_module/add_46/n222 ), .O(\test_module/n1156 [112]), 
            .CO(\test_module/add_46/n224 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i112 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i112 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i113  (.I0(o_pllBr1_reg[113]), .I1(1'b0), 
            .CI(\test_module/add_46/n224 ), .O(\test_module/n1156 [113]), 
            .CO(\test_module/add_46/n226 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i113 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i113 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i114  (.I0(o_pllBr1_reg[114]), .I1(1'b0), 
            .CI(\test_module/add_46/n226 ), .O(\test_module/n1156 [114]), 
            .CO(\test_module/add_46/n228 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i114 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i114 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i115  (.I0(o_pllBr1_reg[115]), .I1(1'b0), 
            .CI(\test_module/add_46/n228 ), .O(\test_module/n1156 [115]), 
            .CO(\test_module/add_46/n230 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i115 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i115 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i116  (.I0(o_pllBr1_reg[116]), .I1(1'b0), 
            .CI(\test_module/add_46/n230 ), .O(\test_module/n1156 [116]), 
            .CO(\test_module/add_46/n232 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i116 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i116 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i117  (.I0(o_pllBr1_reg[117]), .I1(1'b0), 
            .CI(\test_module/add_46/n232 ), .O(\test_module/n1156 [117]), 
            .CO(\test_module/add_46/n234 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i117 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i117 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i118  (.I0(o_pllBr1_reg[118]), .I1(1'b0), 
            .CI(\test_module/add_46/n234 ), .O(\test_module/n1156 [118]), 
            .CO(\test_module/add_46/n236 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i118 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i118 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i119  (.I0(o_pllBr1_reg[119]), .I1(1'b0), 
            .CI(\test_module/add_46/n236 ), .O(\test_module/n1156 [119]), 
            .CO(\test_module/add_46/n238 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i119 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i119 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i120  (.I0(o_pllBr1_reg[120]), .I1(1'b0), 
            .CI(\test_module/add_46/n238 ), .O(\test_module/n1156 [120]), 
            .CO(\test_module/add_46/n240 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i120 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i120 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i121  (.I0(o_pllBr1_reg[121]), .I1(1'b0), 
            .CI(\test_module/add_46/n240 ), .O(\test_module/n1156 [121]), 
            .CO(\test_module/add_46/n242 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i121 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i121 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i122  (.I0(o_pllBr1_reg[122]), .I1(1'b0), 
            .CI(\test_module/add_46/n242 ), .O(\test_module/n1156 [122]), 
            .CO(\test_module/add_46/n244 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i122 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i122 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i123  (.I0(o_pllBr1_reg[123]), .I1(1'b0), 
            .CI(\test_module/add_46/n244 ), .O(\test_module/n1156 [123]), 
            .CO(\test_module/add_46/n246 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i123 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i123 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i124  (.I0(o_pllBr1_reg[124]), .I1(1'b0), 
            .CI(\test_module/add_46/n246 ), .O(\test_module/n1156 [124]), 
            .CO(\test_module/add_46/n248 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i124 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i124 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i125  (.I0(o_pllBr1_reg[125]), .I1(1'b0), 
            .CI(\test_module/add_46/n248 ), .O(\test_module/n1156 [125]), 
            .CO(\test_module/add_46/n250 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i125 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i125 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i126  (.I0(o_pllBr1_reg[126]), .I1(1'b0), 
            .CI(\test_module/add_46/n250 ), .O(\test_module/n1156 [126]), 
            .CO(\test_module/add_46/n252 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i126 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i126 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i127  (.I0(o_pllBr1_reg[127]), .I1(1'b0), 
            .CI(\test_module/add_46/n252 ), .O(\test_module/n1156 [127]), 
            .CO(\test_module/add_46/n254 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i127 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i127 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i128  (.I0(o_pllBr1_reg[128]), .I1(1'b0), 
            .CI(\test_module/add_46/n254 ), .O(\test_module/n1156 [128]), 
            .CO(\test_module/add_46/n256 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i128 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i128 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i129  (.I0(o_pllBr1_reg[129]), .I1(1'b0), 
            .CI(\test_module/add_46/n256 ), .O(\test_module/n1156 [129]), 
            .CO(\test_module/add_46/n258 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i129 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i129 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i130  (.I0(o_pllBr1_reg[130]), .I1(1'b0), 
            .CI(\test_module/add_46/n258 ), .O(\test_module/n1156 [130]), 
            .CO(\test_module/add_46/n260 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i130 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i130 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i131  (.I0(o_pllBr1_reg[131]), .I1(1'b0), 
            .CI(\test_module/add_46/n260 ), .O(\test_module/n1156 [131]), 
            .CO(\test_module/add_46/n262 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i131 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i131 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i132  (.I0(o_pllBr1_reg[132]), .I1(1'b0), 
            .CI(\test_module/add_46/n262 ), .O(\test_module/n1156 [132]), 
            .CO(\test_module/add_46/n264 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i132 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i132 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i133  (.I0(o_pllBr1_reg[133]), .I1(1'b0), 
            .CI(\test_module/add_46/n264 ), .O(\test_module/n1156 [133]), 
            .CO(\test_module/add_46/n266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i133 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i133 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i134  (.I0(o_pllBr1_reg[134]), .I1(1'b0), 
            .CI(\test_module/add_46/n266 ), .O(\test_module/n1156 [134]), 
            .CO(\test_module/add_46/n268 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i134 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i134 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i135  (.I0(o_pllBr1_reg[135]), .I1(1'b0), 
            .CI(\test_module/add_46/n268 ), .O(\test_module/n1156 [135]), 
            .CO(\test_module/add_46/n270 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i135 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i135 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i136  (.I0(o_pllBr1_reg[136]), .I1(1'b0), 
            .CI(\test_module/add_46/n270 ), .O(\test_module/n1156 [136]), 
            .CO(\test_module/add_46/n272 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i136 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i136 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i137  (.I0(o_pllBr1_reg[137]), .I1(1'b0), 
            .CI(\test_module/add_46/n272 ), .O(\test_module/n1156 [137]), 
            .CO(\test_module/add_46/n274 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i137 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i137 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i138  (.I0(o_pllBr1_reg[138]), .I1(1'b0), 
            .CI(\test_module/add_46/n274 ), .O(\test_module/n1156 [138]), 
            .CO(\test_module/add_46/n276 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i138 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i138 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i139  (.I0(o_pllBr1_reg[139]), .I1(1'b0), 
            .CI(\test_module/add_46/n276 ), .O(\test_module/n1156 [139]), 
            .CO(\test_module/add_46/n278 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i139 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i139 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i140  (.I0(o_pllBr1_reg[140]), .I1(1'b0), 
            .CI(\test_module/add_46/n278 ), .O(\test_module/n1156 [140]), 
            .CO(\test_module/add_46/n280 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i140 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i140 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i141  (.I0(o_pllBr1_reg[141]), .I1(1'b0), 
            .CI(\test_module/add_46/n280 ), .O(\test_module/n1156 [141]), 
            .CO(\test_module/add_46/n282 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i141 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i141 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i142  (.I0(o_pllBr1_reg[142]), .I1(1'b0), 
            .CI(\test_module/add_46/n282 ), .O(\test_module/n1156 [142]), 
            .CO(\test_module/add_46/n284 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i142 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i142 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i143  (.I0(o_pllBr1_reg[143]), .I1(1'b0), 
            .CI(\test_module/add_46/n284 ), .O(\test_module/n1156 [143]), 
            .CO(\test_module/add_46/n286 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i143 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i143 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i144  (.I0(o_pllBr1_reg[144]), .I1(1'b0), 
            .CI(\test_module/add_46/n286 ), .O(\test_module/n1156 [144]), 
            .CO(\test_module/add_46/n288 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i144 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i144 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i145  (.I0(o_pllBr1_reg[145]), .I1(1'b0), 
            .CI(\test_module/add_46/n288 ), .O(\test_module/n1156 [145]), 
            .CO(\test_module/add_46/n290 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i145 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i145 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i146  (.I0(o_pllBr1_reg[146]), .I1(1'b0), 
            .CI(\test_module/add_46/n290 ), .O(\test_module/n1156 [146]), 
            .CO(\test_module/add_46/n292 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i146 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i146 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i147  (.I0(o_pllBr1_reg[147]), .I1(1'b0), 
            .CI(\test_module/add_46/n292 ), .O(\test_module/n1156 [147]), 
            .CO(\test_module/add_46/n294 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i147 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i147 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i148  (.I0(o_pllBr1_reg[148]), .I1(1'b0), 
            .CI(\test_module/add_46/n294 ), .O(\test_module/n1156 [148]), 
            .CO(\test_module/add_46/n296 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i148 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i148 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i149  (.I0(o_pllBr1_reg[149]), .I1(1'b0), 
            .CI(\test_module/add_46/n296 ), .O(\test_module/n1156 [149]), 
            .CO(\test_module/add_46/n298 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i149 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i149 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i150  (.I0(o_pllBr1_reg[150]), .I1(1'b0), 
            .CI(\test_module/add_46/n298 ), .O(\test_module/n1156 [150]), 
            .CO(\test_module/add_46/n300 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i150 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i150 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i151  (.I0(o_pllBr1_reg[151]), .I1(1'b0), 
            .CI(\test_module/add_46/n300 ), .O(\test_module/n1156 [151]), 
            .CO(\test_module/add_46/n302 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i151 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i151 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i152  (.I0(o_pllBr1_reg[152]), .I1(1'b0), 
            .CI(\test_module/add_46/n302 ), .O(\test_module/n1156 [152]), 
            .CO(\test_module/add_46/n304 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i152 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i152 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i153  (.I0(o_pllBr1_reg[153]), .I1(1'b0), 
            .CI(\test_module/add_46/n304 ), .O(\test_module/n1156 [153]), 
            .CO(\test_module/add_46/n306 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i153 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i153 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i154  (.I0(o_pllBr1_reg[154]), .I1(1'b0), 
            .CI(\test_module/add_46/n306 ), .O(\test_module/n1156 [154]), 
            .CO(\test_module/add_46/n308 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i154 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i154 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i155  (.I0(o_pllBr1_reg[155]), .I1(1'b0), 
            .CI(\test_module/add_46/n308 ), .O(\test_module/n1156 [155]), 
            .CO(\test_module/add_46/n310 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i155 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i155 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i156  (.I0(o_pllBr1_reg[156]), .I1(1'b0), 
            .CI(\test_module/add_46/n310 ), .O(\test_module/n1156 [156]), 
            .CO(\test_module/add_46/n312 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i156 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i156 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i157  (.I0(o_pllBr1_reg[157]), .I1(1'b0), 
            .CI(\test_module/add_46/n312 ), .O(\test_module/n1156 [157]), 
            .CO(\test_module/add_46/n314 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i157 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i157 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i158  (.I0(o_pllBr1_reg[158]), .I1(1'b0), 
            .CI(\test_module/add_46/n314 ), .O(\test_module/n1156 [158]), 
            .CO(\test_module/add_46/n316 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i158 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i158 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i159  (.I0(o_pllBr1_reg[159]), .I1(1'b0), 
            .CI(\test_module/add_46/n316 ), .O(\test_module/n1156 [159]), 
            .CO(\test_module/add_46/n318 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i159 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i159 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i160  (.I0(o_pllBr1_reg[160]), .I1(1'b0), 
            .CI(\test_module/add_46/n318 ), .O(\test_module/n1156 [160]), 
            .CO(\test_module/add_46/n320 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i160 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i160 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i161  (.I0(o_pllBr1_reg[161]), .I1(1'b0), 
            .CI(\test_module/add_46/n320 ), .O(\test_module/n1156 [161]), 
            .CO(\test_module/add_46/n322 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i161 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i161 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i162  (.I0(o_pllBr1_reg[162]), .I1(1'b0), 
            .CI(\test_module/add_46/n322 ), .O(\test_module/n1156 [162]), 
            .CO(\test_module/add_46/n324 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i162 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i162 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i163  (.I0(o_pllBr1_reg[163]), .I1(1'b0), 
            .CI(\test_module/add_46/n324 ), .O(\test_module/n1156 [163]), 
            .CO(\test_module/add_46/n326 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i163 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i163 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i164  (.I0(o_pllBr1_reg[164]), .I1(1'b0), 
            .CI(\test_module/add_46/n326 ), .O(\test_module/n1156 [164]), 
            .CO(\test_module/add_46/n328 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i164 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i164 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i165  (.I0(o_pllBr1_reg[165]), .I1(1'b0), 
            .CI(\test_module/add_46/n328 ), .O(\test_module/n1156 [165]), 
            .CO(\test_module/add_46/n330 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i165 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i165 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i166  (.I0(o_pllBr1_reg[166]), .I1(1'b0), 
            .CI(\test_module/add_46/n330 ), .O(\test_module/n1156 [166]), 
            .CO(\test_module/add_46/n332 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i166 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i166 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i167  (.I0(o_pllBr1_reg[167]), .I1(1'b0), 
            .CI(\test_module/add_46/n332 ), .O(\test_module/n1156 [167]), 
            .CO(\test_module/add_46/n334 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i167 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i167 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i168  (.I0(o_pllBr1_reg[168]), .I1(1'b0), 
            .CI(\test_module/add_46/n334 ), .O(\test_module/n1156 [168]), 
            .CO(\test_module/add_46/n336 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i168 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i168 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i169  (.I0(o_pllBr1_reg[169]), .I1(1'b0), 
            .CI(\test_module/add_46/n336 ), .O(\test_module/n1156 [169]), 
            .CO(\test_module/add_46/n338 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i169 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i169 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i170  (.I0(o_pllBr1_reg[170]), .I1(1'b0), 
            .CI(\test_module/add_46/n338 ), .O(\test_module/n1156 [170]), 
            .CO(\test_module/add_46/n340 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i170 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i170 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i171  (.I0(o_pllBr1_reg[171]), .I1(1'b0), 
            .CI(\test_module/add_46/n340 ), .O(\test_module/n1156 [171]), 
            .CO(\test_module/add_46/n342 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i171 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i171 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i172  (.I0(o_pllBr1_reg[172]), .I1(1'b0), 
            .CI(\test_module/add_46/n342 ), .O(\test_module/n1156 [172]), 
            .CO(\test_module/add_46/n344 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i172 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i172 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i173  (.I0(o_pllBr1_reg[173]), .I1(1'b0), 
            .CI(\test_module/add_46/n344 ), .O(\test_module/n1156 [173]), 
            .CO(\test_module/add_46/n346 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i173 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i173 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i174  (.I0(o_pllBr1_reg[174]), .I1(1'b0), 
            .CI(\test_module/add_46/n346 ), .O(\test_module/n1156 [174]), 
            .CO(\test_module/add_46/n348 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i174 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i174 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i175  (.I0(o_pllBr1_reg[175]), .I1(1'b0), 
            .CI(\test_module/add_46/n348 ), .O(\test_module/n1156 [175]), 
            .CO(\test_module/add_46/n350 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i175 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i175 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i176  (.I0(o_pllBr1_reg[176]), .I1(1'b0), 
            .CI(\test_module/add_46/n350 ), .O(\test_module/n1156 [176]), 
            .CO(\test_module/add_46/n352 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i176 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i176 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i177  (.I0(o_pllBr1_reg[177]), .I1(1'b0), 
            .CI(\test_module/add_46/n352 ), .O(\test_module/n1156 [177]), 
            .CO(\test_module/add_46/n354 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i177 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i177 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i178  (.I0(o_pllBr1_reg[178]), .I1(1'b0), 
            .CI(\test_module/add_46/n354 ), .O(\test_module/n1156 [178]), 
            .CO(\test_module/add_46/n356 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i178 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i178 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i179  (.I0(o_pllBr1_reg[179]), .I1(1'b0), 
            .CI(\test_module/add_46/n356 ), .O(\test_module/n1156 [179]), 
            .CO(\test_module/add_46/n358 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i179 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i179 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i180  (.I0(o_pllBr1_reg[180]), .I1(1'b0), 
            .CI(\test_module/add_46/n358 ), .O(\test_module/n1156 [180]), 
            .CO(\test_module/add_46/n360 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i180 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i180 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i181  (.I0(o_pllBr1_reg[181]), .I1(1'b0), 
            .CI(\test_module/add_46/n360 ), .O(\test_module/n1156 [181]), 
            .CO(\test_module/add_46/n362 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i181 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i181 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i182  (.I0(o_pllBr1_reg[182]), .I1(1'b0), 
            .CI(\test_module/add_46/n362 ), .O(\test_module/n1156 [182]), 
            .CO(\test_module/add_46/n364 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i182 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i182 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i183  (.I0(o_pllBr1_reg[183]), .I1(1'b0), 
            .CI(\test_module/add_46/n364 ), .O(\test_module/n1156 [183]), 
            .CO(\test_module/add_46/n366 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i183 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i183 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i184  (.I0(o_pllBr1_reg[184]), .I1(1'b0), 
            .CI(\test_module/add_46/n366 ), .O(\test_module/n1156 [184]), 
            .CO(\test_module/add_46/n368 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i184 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i184 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i185  (.I0(o_pllBr1_reg[185]), .I1(1'b0), 
            .CI(\test_module/add_46/n368 ), .O(\test_module/n1156 [185]), 
            .CO(\test_module/add_46/n370 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i185 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i185 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i186  (.I0(o_pllBr1_reg[186]), .I1(1'b0), 
            .CI(\test_module/add_46/n370 ), .O(\test_module/n1156 [186]), 
            .CO(\test_module/add_46/n372 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i186 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i186 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i187  (.I0(o_pllBr1_reg[187]), .I1(1'b0), 
            .CI(\test_module/add_46/n372 ), .O(\test_module/n1156 [187]), 
            .CO(\test_module/add_46/n374 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i187 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i187 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i188  (.I0(o_pllBr1_reg[188]), .I1(1'b0), 
            .CI(\test_module/add_46/n374 ), .O(\test_module/n1156 [188]), 
            .CO(\test_module/add_46/n376 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i188 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i188 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i189  (.I0(o_pllBr1_reg[189]), .I1(1'b0), 
            .CI(\test_module/add_46/n376 ), .O(\test_module/n1156 [189]), 
            .CO(\test_module/add_46/n378 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i189 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i189 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i190  (.I0(o_pllBr1_reg[190]), .I1(1'b0), 
            .CI(\test_module/add_46/n378 ), .O(\test_module/n1156 [190]), 
            .CO(\test_module/add_46/n380 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i190 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i190 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i191  (.I0(o_pllBr1_reg[191]), .I1(1'b0), 
            .CI(\test_module/add_46/n380 ), .O(\test_module/n1156 [191]), 
            .CO(\test_module/add_46/n382 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i191 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i191 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i192  (.I0(o_pllBr1_reg[192]), .I1(1'b0), 
            .CI(\test_module/add_46/n382 ), .O(\test_module/n1156 [192]), 
            .CO(\test_module/add_46/n384 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i192 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i192 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i193  (.I0(o_pllBr1_reg[193]), .I1(1'b0), 
            .CI(\test_module/add_46/n384 ), .O(\test_module/n1156 [193]), 
            .CO(\test_module/add_46/n386 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i193 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i193 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i194  (.I0(o_pllBr1_reg[194]), .I1(1'b0), 
            .CI(\test_module/add_46/n386 ), .O(\test_module/n1156 [194]), 
            .CO(\test_module/add_46/n388 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i194 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i194 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i195  (.I0(o_pllBr1_reg[195]), .I1(1'b0), 
            .CI(\test_module/add_46/n388 ), .O(\test_module/n1156 [195]), 
            .CO(\test_module/add_46/n390 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i195 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i195 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i196  (.I0(o_pllBr1_reg[196]), .I1(1'b0), 
            .CI(\test_module/add_46/n390 ), .O(\test_module/n1156 [196]), 
            .CO(\test_module/add_46/n392 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i196 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i196 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i197  (.I0(o_pllBr1_reg[197]), .I1(1'b0), 
            .CI(\test_module/add_46/n392 ), .O(\test_module/n1156 [197]), 
            .CO(\test_module/add_46/n394 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i197 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i197 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i198  (.I0(o_pllBr1_reg[198]), .I1(1'b0), 
            .CI(\test_module/add_46/n394 ), .O(\test_module/n1156 [198]), 
            .CO(\test_module/add_46/n396 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i198 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i198 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i199  (.I0(o_pllBr1_reg[199]), .I1(1'b0), 
            .CI(\test_module/add_46/n396 ), .O(\test_module/n1156 [199]), 
            .CO(\test_module/add_46/n398 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i199 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i199 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i200  (.I0(o_pllBr1_reg[200]), .I1(1'b0), 
            .CI(\test_module/add_46/n398 ), .O(\test_module/n1156 [200]), 
            .CO(\test_module/add_46/n400 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i200 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i200 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i201  (.I0(o_pllBr1_reg[201]), .I1(1'b0), 
            .CI(\test_module/add_46/n400 ), .O(\test_module/n1156 [201]), 
            .CO(\test_module/add_46/n402 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i201 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i201 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i202  (.I0(o_pllBr1_reg[202]), .I1(1'b0), 
            .CI(\test_module/add_46/n402 ), .O(\test_module/n1156 [202]), 
            .CO(\test_module/add_46/n404 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i202 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i202 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i203  (.I0(o_pllBr1_reg[203]), .I1(1'b0), 
            .CI(\test_module/add_46/n404 ), .O(\test_module/n1156 [203]), 
            .CO(\test_module/add_46/n406 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i203 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i203 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i204  (.I0(o_pllBr1_reg[204]), .I1(1'b0), 
            .CI(\test_module/add_46/n406 ), .O(\test_module/n1156 [204]), 
            .CO(\test_module/add_46/n408 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i204 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i204 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i205  (.I0(o_pllBr1_reg[205]), .I1(1'b0), 
            .CI(\test_module/add_46/n408 ), .O(\test_module/n1156 [205]), 
            .CO(\test_module/add_46/n410 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i205 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i205 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i206  (.I0(o_pllBr1_reg[206]), .I1(1'b0), 
            .CI(\test_module/add_46/n410 ), .O(\test_module/n1156 [206]), 
            .CO(\test_module/add_46/n412 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i206 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i206 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i207  (.I0(o_pllBr1_reg[207]), .I1(1'b0), 
            .CI(\test_module/add_46/n412 ), .O(\test_module/n1156 [207]), 
            .CO(\test_module/add_46/n414 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i207 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i207 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i208  (.I0(o_pllBr1_reg[208]), .I1(1'b0), 
            .CI(\test_module/add_46/n414 ), .O(\test_module/n1156 [208]), 
            .CO(\test_module/add_46/n416 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i208 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i208 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i209  (.I0(o_pllBr1_reg[209]), .I1(1'b0), 
            .CI(\test_module/add_46/n416 ), .O(\test_module/n1156 [209]), 
            .CO(\test_module/add_46/n418 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i209 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i209 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i210  (.I0(o_pllBr1_reg[210]), .I1(1'b0), 
            .CI(\test_module/add_46/n418 ), .O(\test_module/n1156 [210]), 
            .CO(\test_module/add_46/n420 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i210 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i210 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i211  (.I0(o_pllBr1_reg[211]), .I1(1'b0), 
            .CI(\test_module/add_46/n420 ), .O(\test_module/n1156 [211]), 
            .CO(\test_module/add_46/n422 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i211 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i211 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i212  (.I0(o_pllBr1_reg[212]), .I1(1'b0), 
            .CI(\test_module/add_46/n422 ), .O(\test_module/n1156 [212]), 
            .CO(\test_module/add_46/n424 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i212 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i212 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i213  (.I0(o_pllBr1_reg[213]), .I1(1'b0), 
            .CI(\test_module/add_46/n424 ), .O(\test_module/n1156 [213]), 
            .CO(\test_module/add_46/n426 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i213 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i213 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i214  (.I0(o_pllBr1_reg[214]), .I1(1'b0), 
            .CI(\test_module/add_46/n426 ), .O(\test_module/n1156 [214]), 
            .CO(\test_module/add_46/n428 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i214 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i214 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i215  (.I0(o_pllBr1_reg[215]), .I1(1'b0), 
            .CI(\test_module/add_46/n428 ), .O(\test_module/n1156 [215]), 
            .CO(\test_module/add_46/n430 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i215 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i215 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i216  (.I0(o_pllBr1_reg[216]), .I1(1'b0), 
            .CI(\test_module/add_46/n430 ), .O(\test_module/n1156 [216]), 
            .CO(\test_module/add_46/n432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i216 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i216 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i217  (.I0(o_pllBr1_reg[217]), .I1(1'b0), 
            .CI(\test_module/add_46/n432 ), .O(\test_module/n1156 [217]), 
            .CO(\test_module/add_46/n434 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i217 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i217 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i218  (.I0(o_pllBr1_reg[218]), .I1(1'b0), 
            .CI(\test_module/add_46/n434 ), .O(\test_module/n1156 [218]), 
            .CO(\test_module/add_46/n436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i218 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i218 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i219  (.I0(o_pllBr1_reg[219]), .I1(1'b0), 
            .CI(\test_module/add_46/n436 ), .O(\test_module/n1156 [219]), 
            .CO(\test_module/add_46/n438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i219 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i219 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i220  (.I0(o_pllBr1_reg[220]), .I1(1'b0), 
            .CI(\test_module/add_46/n438 ), .O(\test_module/n1156 [220]), 
            .CO(\test_module/add_46/n440 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i220 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i220 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i221  (.I0(o_pllBr1_reg[221]), .I1(1'b0), 
            .CI(\test_module/add_46/n440 ), .O(\test_module/n1156 [221]), 
            .CO(\test_module/add_46/n442 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i221 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i221 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i222  (.I0(o_pllBr1_reg[222]), .I1(1'b0), 
            .CI(\test_module/add_46/n442 ), .O(\test_module/n1156 [222]), 
            .CO(\test_module/add_46/n444 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i222 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i222 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i223  (.I0(o_pllBr1_reg[223]), .I1(1'b0), 
            .CI(\test_module/add_46/n444 ), .O(\test_module/n1156 [223]), 
            .CO(\test_module/add_46/n446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i223 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i223 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i224  (.I0(o_pllBr1_reg[224]), .I1(1'b0), 
            .CI(\test_module/add_46/n446 ), .O(\test_module/n1156 [224]), 
            .CO(\test_module/add_46/n448 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i224 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i224 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i225  (.I0(o_pllBr1_reg[225]), .I1(1'b0), 
            .CI(\test_module/add_46/n448 ), .O(\test_module/n1156 [225]), 
            .CO(\test_module/add_46/n450 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i225 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i225 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i226  (.I0(o_pllBr1_reg[226]), .I1(1'b0), 
            .CI(\test_module/add_46/n450 ), .O(\test_module/n1156 [226]), 
            .CO(\test_module/add_46/n452 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i226 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i226 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i227  (.I0(o_pllBr1_reg[227]), .I1(1'b0), 
            .CI(\test_module/add_46/n452 ), .O(\test_module/n1156 [227]), 
            .CO(\test_module/add_46/n454 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i227 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i227 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i228  (.I0(o_pllBr1_reg[228]), .I1(1'b0), 
            .CI(\test_module/add_46/n454 ), .O(\test_module/n1156 [228]), 
            .CO(\test_module/add_46/n456 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i228 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i228 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i229  (.I0(o_pllBr1_reg[229]), .I1(1'b0), 
            .CI(\test_module/add_46/n456 ), .O(\test_module/n1156 [229]), 
            .CO(\test_module/add_46/n458 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i229 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i229 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i230  (.I0(o_pllBr1_reg[230]), .I1(1'b0), 
            .CI(\test_module/add_46/n458 ), .O(\test_module/n1156 [230]), 
            .CO(\test_module/add_46/n460 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i230 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i230 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i231  (.I0(o_pllBr1_reg[231]), .I1(1'b0), 
            .CI(\test_module/add_46/n460 ), .O(\test_module/n1156 [231]), 
            .CO(\test_module/add_46/n462 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i231 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i231 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i232  (.I0(o_pllBr1_reg[232]), .I1(1'b0), 
            .CI(\test_module/add_46/n462 ), .O(\test_module/n1156 [232]), 
            .CO(\test_module/add_46/n464 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i232 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i232 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i233  (.I0(o_pllBr1_reg[233]), .I1(1'b0), 
            .CI(\test_module/add_46/n464 ), .O(\test_module/n1156 [233]), 
            .CO(\test_module/add_46/n466 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i233 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i233 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i234  (.I0(o_pllBr1_reg[234]), .I1(1'b0), 
            .CI(\test_module/add_46/n466 ), .O(\test_module/n1156 [234]), 
            .CO(\test_module/add_46/n468 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i234 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i234 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i235  (.I0(o_pllBr1_reg[235]), .I1(1'b0), 
            .CI(\test_module/add_46/n468 ), .O(\test_module/n1156 [235]), 
            .CO(\test_module/add_46/n470 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i235 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i235 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i236  (.I0(o_pllBr1_reg[236]), .I1(1'b0), 
            .CI(\test_module/add_46/n470 ), .O(\test_module/n1156 [236]), 
            .CO(\test_module/add_46/n472 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i236 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i236 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i237  (.I0(o_pllBr1_reg[237]), .I1(1'b0), 
            .CI(\test_module/add_46/n472 ), .O(\test_module/n1156 [237]), 
            .CO(\test_module/add_46/n474 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i237 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i237 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i238  (.I0(o_pllBr1_reg[238]), .I1(1'b0), 
            .CI(\test_module/add_46/n474 ), .O(\test_module/n1156 [238]), 
            .CO(\test_module/add_46/n476 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i238 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i238 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i239  (.I0(o_pllBr1_reg[239]), .I1(1'b0), 
            .CI(\test_module/add_46/n476 ), .O(\test_module/n1156 [239]), 
            .CO(\test_module/add_46/n478 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i239 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i239 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i240  (.I0(o_pllBr1_reg[240]), .I1(1'b0), 
            .CI(\test_module/add_46/n478 ), .O(\test_module/n1156 [240]), 
            .CO(\test_module/add_46/n480 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i240 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i240 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i241  (.I0(o_pllBr1_reg[241]), .I1(1'b0), 
            .CI(\test_module/add_46/n480 ), .O(\test_module/n1156 [241]), 
            .CO(\test_module/add_46/n482 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i241 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i241 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i242  (.I0(o_pllBr1_reg[242]), .I1(1'b0), 
            .CI(\test_module/add_46/n482 ), .O(\test_module/n1156 [242]), 
            .CO(\test_module/add_46/n484 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i242 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i242 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i243  (.I0(o_pllBr1_reg[243]), .I1(1'b0), 
            .CI(\test_module/add_46/n484 ), .O(\test_module/n1156 [243]), 
            .CO(\test_module/add_46/n486 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i243 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i243 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i244  (.I0(o_pllBr1_reg[244]), .I1(1'b0), 
            .CI(\test_module/add_46/n486 ), .O(\test_module/n1156 [244]), 
            .CO(\test_module/add_46/n488 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i244 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i244 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i245  (.I0(o_pllBr1_reg[245]), .I1(1'b0), 
            .CI(\test_module/add_46/n488 ), .O(\test_module/n1156 [245]), 
            .CO(\test_module/add_46/n490 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i245 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i245 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i246  (.I0(o_pllBr1_reg[246]), .I1(1'b0), 
            .CI(\test_module/add_46/n490 ), .O(\test_module/n1156 [246]), 
            .CO(\test_module/add_46/n492 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i246 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i246 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i247  (.I0(o_pllBr1_reg[247]), .I1(1'b0), 
            .CI(\test_module/add_46/n492 ), .O(\test_module/n1156 [247]), 
            .CO(\test_module/add_46/n494 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i247 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i247 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i248  (.I0(o_pllBr1_reg[248]), .I1(1'b0), 
            .CI(\test_module/add_46/n494 ), .O(\test_module/n1156 [248]), 
            .CO(\test_module/add_46/n496 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i248 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i248 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i249  (.I0(o_pllBr1_reg[249]), .I1(1'b0), 
            .CI(\test_module/add_46/n496 ), .O(\test_module/n1156 [249]), 
            .CO(\test_module/add_46/n498 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i249 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i249 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i250  (.I0(o_pllBr1_reg[250]), .I1(1'b0), 
            .CI(\test_module/add_46/n498 ), .O(\test_module/n1156 [250]), 
            .CO(\test_module/add_46/n500 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i250 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i250 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i251  (.I0(o_pllBr1_reg[251]), .I1(1'b0), 
            .CI(\test_module/add_46/n500 ), .O(\test_module/n1156 [251]), 
            .CO(\test_module/add_46/n502 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i251 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i251 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i252  (.I0(o_pllBr1_reg[252]), .I1(1'b0), 
            .CI(\test_module/add_46/n502 ), .O(\test_module/n1156 [252]), 
            .CO(\test_module/add_46/n504 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i252 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i252 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i253  (.I0(o_pllBr1_reg[253]), .I1(1'b0), 
            .CI(\test_module/add_46/n504 ), .O(\test_module/n1156 [253]), 
            .CO(\test_module/add_46/n506 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i253 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i253 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i254  (.I0(o_pllBr1_reg[254]), .I1(1'b0), 
            .CI(\test_module/add_46/n506 ), .O(\test_module/n1156 [254]), 
            .CO(\test_module/add_46/n508 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i254 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i254 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_46/i255  (.I0(o_pllBr1_reg[255]), .I1(1'b0), 
            .CI(\test_module/add_46/n508 ), .O(\test_module/n1156 [255])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(36)
    defparam \test_module/add_46/i255 .I0_POLARITY = 1'b1;
    defparam \test_module/add_46/i255 .I1_POLARITY = 1'b1;
    EFX_ADD \debug_inst/vio0/vio_core_inst/add_772/i2  (.I0(\debug_inst/vio0/vio_core_inst/bit_count [2]), 
            .I1(1'b0), .CI(\debug_inst/vio0/vio_core_inst/add_772/n2 ), 
            .O(\debug_inst/vio0/vio_core_inst/n408 [2]), .CO(\debug_inst/vio0/vio_core_inst/add_772/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1429)
    defparam \debug_inst/vio0/vio_core_inst/add_772/i2 .I0_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/add_772/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \debug_inst/vio0/vio_core_inst/add_772/i3  (.I0(\debug_inst/vio0/vio_core_inst/bit_count [3]), 
            .I1(1'b0), .CI(\debug_inst/vio0/vio_core_inst/add_772/n4 ), 
            .O(\debug_inst/vio0/vio_core_inst/n408 [3]), .CO(\debug_inst/vio0/vio_core_inst/add_772/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1429)
    defparam \debug_inst/vio0/vio_core_inst/add_772/i3 .I0_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/add_772/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \debug_inst/vio0/vio_core_inst/add_772/i4  (.I0(\debug_inst/vio0/vio_core_inst/bit_count [4]), 
            .I1(1'b0), .CI(\debug_inst/vio0/vio_core_inst/add_772/n6 ), 
            .O(\debug_inst/vio0/vio_core_inst/n408 [4]), .CO(\debug_inst/vio0/vio_core_inst/add_772/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1429)
    defparam \debug_inst/vio0/vio_core_inst/add_772/i4 .I0_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/add_772/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \debug_inst/vio0/vio_core_inst/add_772/i5  (.I0(\debug_inst/vio0/vio_core_inst/bit_count [5]), 
            .I1(1'b0), .CI(\debug_inst/vio0/vio_core_inst/add_772/n8 ), 
            .O(\debug_inst/vio0/vio_core_inst/n408 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1429)
    defparam \debug_inst/vio0/vio_core_inst/add_772/i5 .I0_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/add_772/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \debug_inst/vio0/vio_core_inst/add_33/i3  (.I0(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I1(1'b0), .CI(\debug_inst/vio0/vio_core_inst/add_33/n4 ), .O(\debug_inst/vio0/vio_core_inst/incremented_address [2]), 
            .CO(\debug_inst/vio0/vio_core_inst/add_33/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1402)
    defparam \debug_inst/vio0/vio_core_inst/add_33/i3 .I0_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/add_33/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \debug_inst/vio0/vio_core_inst/add_33/i4  (.I0(\debug_inst/vio0/vio_core_inst/address_counter [3]), 
            .I1(1'b0), .CI(\debug_inst/vio0/vio_core_inst/add_33/n6 ), .O(\debug_inst/vio0/vio_core_inst/incremented_address [3]), 
            .CO(\debug_inst/vio0/vio_core_inst/add_33/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1402)
    defparam \debug_inst/vio0/vio_core_inst/add_33/i4 .I0_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/add_33/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \debug_inst/vio0/vio_core_inst/add_33/i5  (.I0(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I1(1'b0), .CI(\debug_inst/vio0/vio_core_inst/add_33/n8 ), .O(\debug_inst/vio0/vio_core_inst/incremented_address [4]), 
            .CO(\debug_inst/vio0/vio_core_inst/add_33/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1402)
    defparam \debug_inst/vio0/vio_core_inst/add_33/i5 .I0_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/add_33/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \debug_inst/vio0/vio_core_inst/add_33/i6  (.I0(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I1(1'b0), .CI(\debug_inst/vio0/vio_core_inst/add_33/n10 ), 
            .O(\debug_inst/vio0/vio_core_inst/incremented_address [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1402)
    defparam \debug_inst/vio0/vio_core_inst/add_33/i6 .I0_POLARITY = 1'b1;
    defparam \debug_inst/vio0/vio_core_inst/add_33/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i50  (.I0(o_pllBr0_reg[50]), .I1(1'b0), 
            .CI(\test_module/add_41/n98 ), .O(\test_module/n33 [50]), .CO(\test_module/add_41/n100 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i50 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i50 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i49  (.I0(o_pllBr0_reg[49]), .I1(1'b0), 
            .CI(\test_module/add_41/n96 ), .O(\test_module/n33 [49]), .CO(\test_module/add_41/n98 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i49 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i49 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i48  (.I0(o_pllBr0_reg[48]), .I1(1'b0), 
            .CI(\test_module/add_41/n94 ), .O(\test_module/n33 [48]), .CO(\test_module/add_41/n96 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i48 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i48 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i47  (.I0(o_pllBr0_reg[47]), .I1(1'b0), 
            .CI(\test_module/add_41/n92 ), .O(\test_module/n33 [47]), .CO(\test_module/add_41/n94 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i47 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i47 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i46  (.I0(o_pllBr0_reg[46]), .I1(1'b0), 
            .CI(\test_module/add_41/n90 ), .O(\test_module/n33 [46]), .CO(\test_module/add_41/n92 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i46 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i46 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i45  (.I0(o_pllBr0_reg[45]), .I1(1'b0), 
            .CI(\test_module/add_41/n88 ), .O(\test_module/n33 [45]), .CO(\test_module/add_41/n90 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i45 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i45 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i44  (.I0(o_pllBr0_reg[44]), .I1(1'b0), 
            .CI(\test_module/add_41/n86 ), .O(\test_module/n33 [44]), .CO(\test_module/add_41/n88 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i44 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i44 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i43  (.I0(o_pllBr0_reg[43]), .I1(1'b0), 
            .CI(\test_module/add_41/n84 ), .O(\test_module/n33 [43]), .CO(\test_module/add_41/n86 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i43 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i43 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i42  (.I0(o_pllBr0_reg[42]), .I1(1'b0), 
            .CI(\test_module/add_41/n82 ), .O(\test_module/n33 [42]), .CO(\test_module/add_41/n84 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i42 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i42 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i41  (.I0(o_pllBr0_reg[41]), .I1(1'b0), 
            .CI(\test_module/add_41/n80 ), .O(\test_module/n33 [41]), .CO(\test_module/add_41/n82 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i41 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i41 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i40  (.I0(o_pllBr0_reg[40]), .I1(1'b0), 
            .CI(\test_module/add_41/n78 ), .O(\test_module/n33 [40]), .CO(\test_module/add_41/n80 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i40 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i40 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i39  (.I0(o_pllBr0_reg[39]), .I1(1'b0), 
            .CI(\test_module/add_41/n76 ), .O(\test_module/n33 [39]), .CO(\test_module/add_41/n78 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i39 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i39 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i87  (.I0(o_pllBr0_reg[87]), .I1(1'b0), 
            .CI(\test_module/add_41/n172 ), .O(\test_module/n33 [87]), .CO(\test_module/add_41/n174 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i87 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i87 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i38  (.I0(o_pllBr0_reg[38]), .I1(1'b0), 
            .CI(\test_module/add_41/n74 ), .O(\test_module/n33 [38]), .CO(\test_module/add_41/n76 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i38 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i38 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i37  (.I0(o_pllBr0_reg[37]), .I1(1'b0), 
            .CI(\test_module/add_41/n72 ), .O(\test_module/n33 [37]), .CO(\test_module/add_41/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i37 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i37 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i36  (.I0(o_pllBr0_reg[36]), .I1(1'b0), 
            .CI(\test_module/add_41/n70 ), .O(\test_module/n33 [36]), .CO(\test_module/add_41/n72 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i36 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i36 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i35  (.I0(o_pllBr0_reg[35]), .I1(1'b0), 
            .CI(\test_module/add_41/n68 ), .O(\test_module/n33 [35]), .CO(\test_module/add_41/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i35 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i35 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i34  (.I0(o_pllBr0_reg[34]), .I1(1'b0), 
            .CI(\test_module/add_41/n66 ), .O(\test_module/n33 [34]), .CO(\test_module/add_41/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i34 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i34 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i33  (.I0(o_pllBr0_reg[33]), .I1(1'b0), 
            .CI(\test_module/add_41/n64 ), .O(\test_module/n33 [33]), .CO(\test_module/add_41/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i33 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i33 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i32  (.I0(o_pllBr0_reg[32]), .I1(1'b0), 
            .CI(\test_module/add_41/n62 ), .O(\test_module/n33 [32]), .CO(\test_module/add_41/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i32 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i31  (.I0(o_pllBr0_reg[31]), .I1(1'b0), 
            .CI(\test_module/add_41/n60 ), .O(\test_module/n33 [31]), .CO(\test_module/add_41/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i31 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i30  (.I0(o_pllBr0_reg[30]), .I1(1'b0), 
            .CI(\test_module/add_41/n58 ), .O(\test_module/n33 [30]), .CO(\test_module/add_41/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i30 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i29  (.I0(o_pllBr0_reg[29]), .I1(1'b0), 
            .CI(\test_module/add_41/n56 ), .O(\test_module/n33 [29]), .CO(\test_module/add_41/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i29 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i28  (.I0(o_pllBr0_reg[28]), .I1(1'b0), 
            .CI(\test_module/add_41/n54 ), .O(\test_module/n33 [28]), .CO(\test_module/add_41/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i28 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i27  (.I0(o_pllBr0_reg[27]), .I1(1'b0), 
            .CI(\test_module/add_41/n52 ), .O(\test_module/n33 [27]), .CO(\test_module/add_41/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i27 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i26  (.I0(o_pllBr0_reg[26]), .I1(1'b0), 
            .CI(\test_module/add_41/n50 ), .O(\test_module/n33 [26]), .CO(\test_module/add_41/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i26 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i25  (.I0(o_pllBr0_reg[25]), .I1(1'b0), 
            .CI(\test_module/add_41/n48 ), .O(\test_module/n33 [25]), .CO(\test_module/add_41/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i25 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i24  (.I0(o_pllBr0_reg[24]), .I1(1'b0), 
            .CI(\test_module/add_41/n46 ), .O(\test_module/n33 [24]), .CO(\test_module/add_41/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i24 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i23  (.I0(o_pllBr0_reg[23]), .I1(1'b0), 
            .CI(\test_module/add_41/n44 ), .O(\test_module/n33 [23]), .CO(\test_module/add_41/n46 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i23 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i22  (.I0(o_pllBr0_reg[22]), .I1(1'b0), 
            .CI(\test_module/add_41/n42 ), .O(\test_module/n33 [22]), .CO(\test_module/add_41/n44 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i22 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i21  (.I0(o_pllBr0_reg[21]), .I1(1'b0), 
            .CI(\test_module/add_41/n40 ), .O(\test_module/n33 [21]), .CO(\test_module/add_41/n42 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i21 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i20  (.I0(o_pllBr0_reg[20]), .I1(1'b0), 
            .CI(\test_module/add_41/n38 ), .O(\test_module/n33 [20]), .CO(\test_module/add_41/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i20 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i19  (.I0(o_pllBr0_reg[19]), .I1(1'b0), 
            .CI(\test_module/add_41/n36 ), .O(\test_module/n33 [19]), .CO(\test_module/add_41/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i19 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i18  (.I0(o_pllBr0_reg[18]), .I1(1'b0), 
            .CI(\test_module/add_41/n34 ), .O(\test_module/n33 [18]), .CO(\test_module/add_41/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i18 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i17  (.I0(o_pllBr0_reg[17]), .I1(1'b0), 
            .CI(\test_module/add_41/n32 ), .O(\test_module/n33 [17]), .CO(\test_module/add_41/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i17 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i16  (.I0(o_pllBr0_reg[16]), .I1(1'b0), 
            .CI(\test_module/add_41/n30 ), .O(\test_module/n33 [16]), .CO(\test_module/add_41/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i16 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i15  (.I0(o_pllBr0_reg[15]), .I1(1'b0), 
            .CI(\test_module/add_41/n28 ), .O(\test_module/n33 [15]), .CO(\test_module/add_41/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i15 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i14  (.I0(o_pllBr0_reg[14]), .I1(1'b0), 
            .CI(\test_module/add_41/n26 ), .O(\test_module/n33 [14]), .CO(\test_module/add_41/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i14 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i13  (.I0(o_pllBr0_reg[13]), .I1(1'b0), 
            .CI(\test_module/add_41/n24 ), .O(\test_module/n33 [13]), .CO(\test_module/add_41/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i13 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i12  (.I0(o_pllBr0_reg[12]), .I1(1'b0), 
            .CI(\test_module/add_41/n22 ), .O(\test_module/n33 [12]), .CO(\test_module/add_41/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i12 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i11  (.I0(o_pllBr0_reg[11]), .I1(1'b0), 
            .CI(\test_module/add_41/n20 ), .O(\test_module/n33 [11]), .CO(\test_module/add_41/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i11 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i10  (.I0(o_pllBr0_reg[10]), .I1(1'b0), 
            .CI(\test_module/add_41/n18 ), .O(\test_module/n33 [10]), .CO(\test_module/add_41/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i10 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i9  (.I0(o_pllBr0_reg[9]), .I1(1'b0), .CI(\test_module/add_41/n16 ), 
            .O(\test_module/n33 [9]), .CO(\test_module/add_41/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i9 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i8  (.I0(o_pllBr0_reg[8]), .I1(1'b0), .CI(\test_module/add_41/n14 ), 
            .O(\test_module/n33 [8]), .CO(\test_module/add_41/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i8 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i7  (.I0(o_pllBr0_reg[7]), .I1(1'b0), .CI(\test_module/add_41/n12 ), 
            .O(\test_module/n33 [7]), .CO(\test_module/add_41/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i7 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i6  (.I0(o_pllBr0_reg[6]), .I1(1'b0), .CI(\test_module/add_41/n10 ), 
            .O(\test_module/n33 [6]), .CO(\test_module/add_41/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i6 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i5  (.I0(o_pllBr0_reg[5]), .I1(1'b0), .CI(\test_module/add_41/n8 ), 
            .O(\test_module/n33 [5]), .CO(\test_module/add_41/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i5 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i4  (.I0(o_pllBr0_reg[4]), .I1(1'b0), .CI(\test_module/add_41/n6 ), 
            .O(\test_module/n33 [4]), .CO(\test_module/add_41/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i4 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i3  (.I0(o_pllBr0_reg[3]), .I1(1'b0), .CI(\test_module/add_41/n4 ), 
            .O(\test_module/n33 [3]), .CO(\test_module/add_41/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i3 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i2  (.I0(o_pllBr0_reg[2]), .I1(1'b0), .CI(\test_module/add_41/n2 ), 
            .O(\test_module/n33 [2]), .CO(\test_module/add_41/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i2 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_39/i13  (.I0(\test_module/delay_1 [13]), .I1(1'b0), 
            .CI(\test_module/add_39/n24 ), .O(\test_module/n9 [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(19)
    defparam \test_module/add_39/i13 .I0_POLARITY = 1'b1;
    defparam \test_module/add_39/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_39/i12  (.I0(\test_module/delay_1 [12]), .I1(1'b0), 
            .CI(\test_module/add_39/n22 ), .O(\test_module/n9 [12]), .CO(\test_module/add_39/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(19)
    defparam \test_module/add_39/i12 .I0_POLARITY = 1'b1;
    defparam \test_module/add_39/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_39/i11  (.I0(\test_module/delay_1 [11]), .I1(1'b0), 
            .CI(\test_module/add_39/n20 ), .O(\test_module/n9 [11]), .CO(\test_module/add_39/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(19)
    defparam \test_module/add_39/i11 .I0_POLARITY = 1'b1;
    defparam \test_module/add_39/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_39/i10  (.I0(\test_module/delay_1 [10]), .I1(1'b0), 
            .CI(\test_module/add_39/n18 ), .O(\test_module/n9 [10]), .CO(\test_module/add_39/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(19)
    defparam \test_module/add_39/i10 .I0_POLARITY = 1'b1;
    defparam \test_module/add_39/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_39/i9  (.I0(\test_module/delay_1 [9]), .I1(1'b0), 
            .CI(\test_module/add_39/n16 ), .O(\test_module/n9 [9]), .CO(\test_module/add_39/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(19)
    defparam \test_module/add_39/i9 .I0_POLARITY = 1'b1;
    defparam \test_module/add_39/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_39/i8  (.I0(\test_module/delay_1 [8]), .I1(1'b0), 
            .CI(\test_module/add_39/n14 ), .O(\test_module/n9 [8]), .CO(\test_module/add_39/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(19)
    defparam \test_module/add_39/i8 .I0_POLARITY = 1'b1;
    defparam \test_module/add_39/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_39/i7  (.I0(\test_module/delay_1 [7]), .I1(1'b0), 
            .CI(\test_module/add_39/n12 ), .O(\test_module/n9 [7]), .CO(\test_module/add_39/n14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(19)
    defparam \test_module/add_39/i7 .I0_POLARITY = 1'b1;
    defparam \test_module/add_39/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_39/i6  (.I0(\test_module/delay_1 [6]), .I1(1'b0), 
            .CI(\test_module/add_39/n10 ), .O(\test_module/n9 [6]), .CO(\test_module/add_39/n12 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(19)
    defparam \test_module/add_39/i6 .I0_POLARITY = 1'b1;
    defparam \test_module/add_39/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_39/i5  (.I0(\test_module/delay_1 [5]), .I1(1'b0), 
            .CI(\test_module/add_39/n8 ), .O(\test_module/n9 [5]), .CO(\test_module/add_39/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(19)
    defparam \test_module/add_39/i5 .I0_POLARITY = 1'b1;
    defparam \test_module/add_39/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_39/i4  (.I0(\test_module/delay_1 [4]), .I1(1'b0), 
            .CI(\test_module/add_39/n6 ), .O(\test_module/n9 [4]), .CO(\test_module/add_39/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(19)
    defparam \test_module/add_39/i4 .I0_POLARITY = 1'b1;
    defparam \test_module/add_39/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_39/i3  (.I0(\test_module/delay_1 [3]), .I1(1'b0), 
            .CI(\test_module/add_39/n4 ), .O(\test_module/n9 [3]), .CO(\test_module/add_39/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(19)
    defparam \test_module/add_39/i3 .I0_POLARITY = 1'b1;
    defparam \test_module/add_39/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_39/i2  (.I0(\test_module/delay_1 [2]), .I1(1'b0), 
            .CI(\test_module/add_39/n2 ), .O(\test_module/n9 [2]), .CO(\test_module/add_39/n4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(19)
    defparam \test_module/add_39/i2 .I0_POLARITY = 1'b1;
    defparam \test_module/add_39/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i94  (.I0(o_pllBr0_reg[94]), .I1(1'b0), 
            .CI(\test_module/add_41/n186 ), .O(\test_module/n33 [94]), .CO(\test_module/add_41/n188 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i94 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i94 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_41/i93  (.I0(o_pllBr0_reg[93]), .I1(1'b0), 
            .CI(\test_module/add_41/n184 ), .O(\test_module/n33 [93]), .CO(\test_module/add_41/n186 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(21)
    defparam \test_module/add_41/i93 .I0_POLARITY = 1'b1;
    defparam \test_module/add_41/i93 .I1_POLARITY = 1'b1;
    EFX_ADD \test_module/add_39/i1  (.I0(\test_module/delay_1 [1]), .I1(\test_module/delay_1 [0]), 
            .CI(1'b0), .O(\test_module/n9 [1]), .CO(\test_module/add_39/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(19)
    defparam \test_module/add_39/i1 .I0_POLARITY = 1'b1;
    defparam \test_module/add_39/i1 .I1_POLARITY = 1'b1;
    EFX_LUT4 LUT__10219 (.I0(\debug_inst/vio0/vio_core_inst/crc_data_out [31]), 
            .I1(\debug_inst/edb_user_dr [81]), .I2(\debug_inst/edb_user_dr [58]), 
            .I3(\debug_inst/vio0/vio_core_inst/crc_data_out [8]), .O(n4095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__10219.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__10220 (.I0(\debug_inst/vio0/vio_core_inst/crc_data_out [22]), 
            .I1(\debug_inst/edb_user_dr [72]), .I2(\debug_inst/edb_user_dr [60]), 
            .I3(\debug_inst/vio0/vio_core_inst/crc_data_out [10]), .O(n4096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__10220.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__10221 (.I0(n4093), .I1(n4094), .I2(n4095), .I3(n4096), 
            .O(n4097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10221.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10222 (.I0(\debug_inst/vio0/vio_core_inst/crc_data_out [25]), 
            .I1(\debug_inst/edb_user_dr [75]), .I2(\debug_inst/edb_user_dr [61]), 
            .I3(\debug_inst/vio0/vio_core_inst/crc_data_out [11]), .O(n4098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__10222.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__10223 (.I0(\debug_inst/vio0/vio_core_inst/crc_data_out [9]), 
            .I1(\debug_inst/edb_user_dr [59]), .I2(\debug_inst/edb_user_dr [52]), 
            .I3(\debug_inst/vio0/vio_core_inst/crc_data_out [2]), .O(n4099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__10223.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__10224 (.I0(\debug_inst/vio0/vio_core_inst/crc_data_out [23]), 
            .I1(\debug_inst/edb_user_dr [73]), .I2(\debug_inst/edb_user_dr [57]), 
            .I3(\debug_inst/vio0/vio_core_inst/crc_data_out [7]), .O(n4100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__10224.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__10225 (.I0(\debug_inst/vio0/vio_core_inst/crc_data_out [6]), 
            .I1(\debug_inst/edb_user_dr [56]), .I2(\debug_inst/edb_user_dr [53]), 
            .I3(\debug_inst/vio0/vio_core_inst/crc_data_out [3]), .O(n4101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__10225.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__10226 (.I0(n4098), .I1(n4099), .I2(n4100), .I3(n4101), 
            .O(n4102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10226.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10227 (.I0(\debug_inst/vio0/vio_core_inst/crc_data_out [26]), 
            .I1(\debug_inst/edb_user_dr [76]), .I2(\debug_inst/edb_user_dr [67]), 
            .I3(\debug_inst/vio0/vio_core_inst/crc_data_out [17]), .O(n4103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__10227.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__10228 (.I0(\debug_inst/vio0/vio_core_inst/crc_data_out [15]), 
            .I1(\debug_inst/edb_user_dr [65]), .I2(\debug_inst/edb_user_dr [64]), 
            .I3(\debug_inst/vio0/vio_core_inst/crc_data_out [14]), .O(n4104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__10228.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__10229 (.I0(\debug_inst/vio0/vio_core_inst/crc_data_out [27]), 
            .I1(\debug_inst/edb_user_dr [77]), .I2(\debug_inst/edb_user_dr [62]), 
            .I3(\debug_inst/vio0/vio_core_inst/crc_data_out [12]), .O(n4105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__10229.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__10230 (.I0(\debug_inst/vio0/vio_core_inst/crc_data_out [30]), 
            .I1(\debug_inst/edb_user_dr [80]), .I2(\debug_inst/edb_user_dr [55]), 
            .I3(\debug_inst/vio0/vio_core_inst/crc_data_out [5]), .O(n4106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__10230.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__10231 (.I0(n4103), .I1(n4104), .I2(n4105), .I3(n4106), 
            .O(n4107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10231.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10232 (.I0(\debug_inst/vio0/vio_core_inst/crc_data_out [16]), 
            .I1(\debug_inst/edb_user_dr [66]), .I2(\debug_inst/edb_user_dr [51]), 
            .I3(\debug_inst/vio0/vio_core_inst/crc_data_out [1]), .O(n4108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__10232.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__10233 (.I0(\debug_inst/vio0/vio_core_inst/crc_data_out [29]), 
            .I1(\debug_inst/edb_user_dr [79]), .I2(\debug_inst/edb_user_dr [71]), 
            .I3(\debug_inst/vio0/vio_core_inst/crc_data_out [21]), .O(n4109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__10233.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__10234 (.I0(\debug_inst/vio0/vio_core_inst/crc_data_out [19]), 
            .I1(\debug_inst/edb_user_dr [69]), .I2(\debug_inst/edb_user_dr [68]), 
            .I3(\debug_inst/vio0/vio_core_inst/crc_data_out [18]), .O(n4110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__10234.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__10235 (.I0(\debug_inst/vio0/vio_core_inst/crc_data_out [13]), 
            .I1(\debug_inst/edb_user_dr [63]), .I2(\debug_inst/edb_user_dr [50]), 
            .I3(\debug_inst/vio0/vio_core_inst/crc_data_out [0]), .O(n4111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__10235.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__10236 (.I0(n4108), .I1(n4109), .I2(n4110), .I3(n4111), 
            .O(n4112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10236.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10237 (.I0(n4097), .I1(n4102), .I2(n4107), .I3(n4112), 
            .O(n4113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10237.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10238 (.I0(\debug_inst/vio0/vio_core_inst/module_state [0]), 
            .I1(\debug_inst/vio0/vio_core_inst/module_state [1]), .O(n4114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10238.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10239 (.I0(\debug_inst/vio0/vio_core_inst/bit_count [0]), 
            .I1(\debug_inst/vio0/vio_core_inst/bit_count [3]), .I2(\debug_inst/vio0/vio_core_inst/bit_count [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/bit_count [1]), .O(n4115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10239.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10240 (.I0(bscan_UPDATE), .I1(\debug_inst/vio0/vio_core_inst/bit_count [4]), 
            .I2(\debug_inst/vio0/vio_core_inst/bit_count [5]), .I3(n4115), 
            .O(n4116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10240.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10241 (.I0(\debug_inst/vio0/vio_core_inst/module_state [1]), 
            .I1(\debug_inst/vio0/vio_core_inst/module_state [3]), .I2(\debug_inst/vio0/vio_core_inst/module_state [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/module_state [0]), .O(n4117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10241.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10242 (.I0(n4116), .I1(n4114), .I2(n4117), .O(n4118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__10242.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__10243 (.I0(n4113), .I1(n4118), .I2(\debug_inst/vio0/vio_core_inst/module_state [3]), 
            .I3(\debug_inst/vio0/vio_core_inst/module_state [1]), .O(n4119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10243.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10244 (.I0(\debug_inst/vio0/vio_core_inst/module_state [2]), 
            .I1(\debug_inst/vio0/vio_core_inst/module_state [3]), .O(n4120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10244.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10245 (.I0(n4120), .I1(\debug_inst/vio0/vio_core_inst/module_state [0]), 
            .O(n4121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10245.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10246 (.I0(\debug_inst/vio0/vio_core_inst/crc_data_out [0]), 
            .I1(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [0]), .I2(n4118), 
            .I3(n4121), .O(n4122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10246.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10247 (.I0(\debug_inst/debug_hub_inst/module_id_reg [1]), 
            .I1(\debug_inst/debug_hub_inst/module_id_reg [2]), .I2(\debug_inst/debug_hub_inst/module_id_reg [3]), 
            .I3(\debug_inst/debug_hub_inst/module_id_reg [0]), .O(n4123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10247.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10248 (.I0(n4119), .I1(n4122), .I2(n4123), .O(bscan_TDO)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(466)
    defparam LUT__10248.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10249 (.I0(\test_module/delay_1 [4]), .I1(\test_module/delay_1 [5]), 
            .I2(\test_module/delay_1 [6]), .I3(\test_module/delay_1 [7]), 
            .O(n4124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10249.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10250 (.I0(\test_module/delay_1 [0]), .I1(\test_module/delay_1 [1]), 
            .I2(\test_module/delay_1 [2]), .I3(\test_module/delay_1 [3]), 
            .O(n4125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10250.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10251 (.I0(\test_module/delay_1 [8]), .I1(\test_module/delay_1 [9]), 
            .I2(\test_module/delay_1 [10]), .O(n4126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10251.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10252 (.I0(n4125), .I1(n4124), .I2(n4126), .O(n4127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__10252.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__10253 (.I0(\test_module/delay_1 [12]), .I1(n4127), .I2(\test_module/delay_1 [11]), 
            .I3(\test_module/delay_1 [13]), .O(n4128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10253.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10254 (.I0(n4128), .I1(\test_module/delay_1 [0]), .O(\test_module/n569 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(23)
    defparam LUT__10254.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__10255 (.I0(\test_module/delay_1 [11]), .I1(\test_module/delay_1 [12]), 
            .I2(n4126), .I3(\test_module/delay_1 [13]), .O(n4129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10255.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10256 (.I0(n4129), .I1(n4125), .I2(n4124), .O(\~test_module/equal_8/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10256.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10257 (.I0(\~test_module/equal_8/n41 ), .I1(n4128), .O(ceg_net2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10257.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10258 (.I0(\test_module/delay_2 [0]), .I1(\test_module/delay_2 [1]), 
            .I2(\test_module/delay_2 [2]), .I3(\test_module/delay_2 [3]), 
            .O(n4130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10258.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10259 (.I0(n4130), .I1(\test_module/delay_2 [8]), .I2(\test_module/delay_2 [9]), 
            .I3(\test_module/delay_2 [10]), .O(n4131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10259.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10260 (.I0(\test_module/delay_2 [4]), .I1(\test_module/delay_2 [5]), 
            .I2(\test_module/delay_2 [6]), .I3(\test_module/delay_2 [7]), 
            .O(n4132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10260.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10261 (.I0(\test_module/delay_2 [11]), .I1(\test_module/delay_2 [12]), 
            .O(n4133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__10261.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__10262 (.I0(n4131), .I1(n4132), .I2(n4133), .I3(\test_module/delay_2 [13]), 
            .O(\~test_module/equal_21/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10262.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10263 (.I0(n4132), .I1(\test_module/delay_2 [8]), .I2(\test_module/delay_2 [9]), 
            .I3(\test_module/delay_2 [10]), .O(n4134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10263.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10264 (.I0(n4131), .I1(n4134), .I2(n4133), .I3(\test_module/delay_2 [13]), 
            .O(n4135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10264.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10265 (.I0(n4135), .I1(\test_module/delay_2 [0]), .O(\test_module/n1692 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(38)
    defparam LUT__10265.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__10266 (.I0(\~test_module/equal_21/n41 ), .I1(n4135), .O(ceg_net5)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10266.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10267 (.I0(n4128), .I1(\test_module/n9 [1]), .O(\test_module/n569 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(23)
    defparam LUT__10267.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10268 (.I0(n4128), .I1(\test_module/n9 [2]), .O(\test_module/n569 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(23)
    defparam LUT__10268.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10269 (.I0(n4128), .I1(\test_module/n9 [3]), .O(\test_module/n569 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(23)
    defparam LUT__10269.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10270 (.I0(n4128), .I1(\test_module/n9 [4]), .O(\test_module/n569 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(23)
    defparam LUT__10270.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10271 (.I0(n4128), .I1(\test_module/n9 [5]), .O(\test_module/n569 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(23)
    defparam LUT__10271.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10272 (.I0(n4128), .I1(\test_module/n9 [6]), .O(\test_module/n569 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(23)
    defparam LUT__10272.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10273 (.I0(n4128), .I1(\test_module/n9 [7]), .O(\test_module/n569 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(23)
    defparam LUT__10273.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10274 (.I0(n4128), .I1(\test_module/n9 [8]), .O(\test_module/n569 [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(23)
    defparam LUT__10274.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10275 (.I0(n4128), .I1(\test_module/n9 [9]), .O(\test_module/n569 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(23)
    defparam LUT__10275.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10276 (.I0(n4128), .I1(\test_module/n9 [10]), .O(\test_module/n569 [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(23)
    defparam LUT__10276.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10277 (.I0(n4128), .I1(\test_module/n9 [11]), .O(\test_module/n569 [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(23)
    defparam LUT__10277.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10278 (.I0(n4128), .I1(\test_module/n9 [12]), .O(\test_module/n569 [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(23)
    defparam LUT__10278.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10279 (.I0(n4128), .I1(\test_module/n9 [13]), .O(\test_module/n569 [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(23)
    defparam LUT__10279.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10280 (.I0(n4135), .I1(\test_module/n1132 [1]), .O(\test_module/n1692 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(38)
    defparam LUT__10280.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10281 (.I0(n4135), .I1(\test_module/n1132 [2]), .O(\test_module/n1692 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(38)
    defparam LUT__10281.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10282 (.I0(n4135), .I1(\test_module/n1132 [3]), .O(\test_module/n1692 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(38)
    defparam LUT__10282.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10283 (.I0(n4135), .I1(\test_module/n1132 [4]), .O(\test_module/n1692 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(38)
    defparam LUT__10283.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10284 (.I0(n4135), .I1(\test_module/n1132 [5]), .O(\test_module/n1692 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(38)
    defparam LUT__10284.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10285 (.I0(n4135), .I1(\test_module/n1132 [6]), .O(\test_module/n1692 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(38)
    defparam LUT__10285.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10286 (.I0(n4135), .I1(\test_module/n1132 [7]), .O(\test_module/n1692 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(38)
    defparam LUT__10286.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10287 (.I0(n4135), .I1(\test_module/n1132 [8]), .O(\test_module/n1692 [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(38)
    defparam LUT__10287.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10288 (.I0(n4135), .I1(\test_module/n1132 [9]), .O(\test_module/n1692 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(38)
    defparam LUT__10288.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10289 (.I0(n4135), .I1(\test_module/n1132 [10]), .O(\test_module/n1692 [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(38)
    defparam LUT__10289.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10290 (.I0(n4135), .I1(\test_module/n1132 [11]), .O(\test_module/n1692 [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(38)
    defparam LUT__10290.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10291 (.I0(n4135), .I1(\test_module/n1132 [12]), .O(\test_module/n1692 [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(38)
    defparam LUT__10291.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10292 (.I0(n4135), .I1(\test_module/n1132 [13]), .O(\test_module/n1692 [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/test_counter.v(38)
    defparam LUT__10292.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10293 (.I0(\debug_inst/edb_user_dr [73]), .I1(\debug_inst/edb_user_dr [74]), 
            .I2(\debug_inst/edb_user_dr [75]), .I3(\debug_inst/edb_user_dr [76]), 
            .O(n4136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10293.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10294 (.I0(\debug_inst/vio0/vio_core_inst/module_state [3]), 
            .I1(\debug_inst/vio0/vio_core_inst/module_state [2]), .O(n4137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__10294.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__10295 (.I0(\debug_inst/vio0/vio_core_inst/module_state [0]), 
            .I1(\debug_inst/vio0/vio_core_inst/module_state [1]), .O(n4138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__10295.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__10296 (.I0(n4137), .I1(n4138), .O(n4139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10296.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10297 (.I0(\debug_inst/edb_user_dr [81]), .I1(n4123), 
            .I2(bscan_UPDATE), .I3(n4139), .O(n4140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10297.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10298 (.I0(\debug_inst/edb_user_dr [78]), .I1(\debug_inst/edb_user_dr [77]), 
            .I2(n4140), .I3(\debug_inst/edb_user_dr [80]), .O(\debug_inst/vio0/vio_core_inst/regsel_ld_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1658)
    defparam LUT__10298.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10299 (.I0(\debug_inst/edb_user_dr [79]), .I1(n4136), 
            .I2(\debug_inst/vio0/vio_core_inst/regsel_ld_en ), .O(\debug_inst/vio0/vio_core_inst/n251 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1393)
    defparam LUT__10299.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10300 (.I0(\debug_inst/vio0/vio_core_inst/bit_count [0]), 
            .I1(\debug_inst/vio0/vio_core_inst/bit_count [3]), .I2(\debug_inst/vio0/vio_core_inst/bit_count [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/bit_count [1]), .O(n4141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10300.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10301 (.I0(\debug_inst/vio0/vio_core_inst/bit_count [5]), 
            .I1(\debug_inst/vio0/vio_core_inst/bit_count [4]), .O(n4142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__10301.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__10302 (.I0(n4115), .I1(n4141), .I2(\debug_inst/vio0/vio_core_inst/opcode [1]), 
            .I3(n4142), .O(n4143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__10302.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__10303 (.I0(\debug_inst/vio0/vio_core_inst/module_state [3]), 
            .I1(\debug_inst/vio0/vio_core_inst/module_state [2]), .O(n4144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10303.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10304 (.I0(\debug_inst/vio0/vio_core_inst/module_state [0]), 
            .I1(\debug_inst/vio0/vio_core_inst/module_state [1]), .I2(n4143), 
            .I3(n4144), .O(n4145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__10304.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__10305 (.I0(\debug_inst/edb_user_dr [79]), .I1(n4138), 
            .O(n4146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10305.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10306 (.I0(\debug_inst/edb_user_dr [77]), .I1(\debug_inst/edb_user_dr [80]), 
            .I2(\debug_inst/edb_user_dr [78]), .I3(bscan_UPDATE), .O(n4147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10306.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10307 (.I0(\debug_inst/edb_user_dr [81]), .I1(n4147), 
            .I2(n4123), .O(n4148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10307.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10308 (.I0(\debug_inst/vio0/vio_core_inst/module_state [0]), 
            .I1(\debug_inst/vio0/vio_core_inst/module_state [1]), .O(n4149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10308.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10309 (.I0(bscan_UPDATE), .I1(n4149), .O(n4150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10309.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10310 (.I0(n4148), .I1(n4146), .I2(n4150), .I3(n4137), 
            .O(n4151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__10310.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__10311 (.I0(n4139), .I1(n4148), .O(n4152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10311.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10312 (.I0(n4120), .I1(n4138), .O(n4153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10312.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10313 (.I0(n4145), .I1(n4151), .I2(n4152), .I3(n4153), 
            .O(n4154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10313.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10314 (.I0(\debug_inst/vio0/vio_core_inst/bit_count [0]), 
            .I1(n4154), .O(\debug_inst/vio0/vio_core_inst/n422 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1429)
    defparam LUT__10314.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10315 (.I0(bscan_UPDATE), .I1(\debug_inst/vio0/vio_core_inst/module_state [0]), 
            .I2(n4123), .I3(\debug_inst/edb_user_dr [81]), .O(n4155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10315.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10316 (.I0(n4155), .I1(\debug_inst/vio0/vio_core_inst/module_state [0]), 
            .I2(\debug_inst/vio0/vio_core_inst/module_state [1]), .I3(n4144), 
            .O(n4156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb00 */ ;
    defparam LUT__10316.LUTMASK = 16'heb00;
    EFX_LUT4 LUT__10317 (.I0(n4120), .I1(\debug_inst/vio0/vio_core_inst/module_state [0]), 
            .I2(n4156), .O(n4157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__10317.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__10318 (.I0(n4157), .I1(bscan_SHIFT), .I2(n4154), .O(ceg_net8)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__10318.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__10320 (.I0(\debug_inst/vio0/vio_core_inst/word_count [0]), 
            .I1(\debug_inst/vio0/vio_core_inst/word_count [3]), .I2(\debug_inst/vio0/vio_core_inst/word_count [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/word_count [1]), .O(n4158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10320.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10321 (.I0(\debug_inst/vio0/vio_core_inst/word_count [7]), 
            .I1(\debug_inst/vio0/vio_core_inst/word_count [6]), .I2(\debug_inst/vio0/vio_core_inst/word_count [5]), 
            .I3(\debug_inst/vio0/vio_core_inst/word_count [4]), .O(n4159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10321.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10322 (.I0(n4158), .I1(n4159), .O(n4160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10322.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10323 (.I0(n4160), .I1(\debug_inst/vio0/vio_core_inst/word_count [8]), 
            .I2(\debug_inst/vio0/vio_core_inst/word_count [9]), .O(n4161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__10323.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__10324 (.I0(\debug_inst/vio0/vio_core_inst/word_count [12]), 
            .I1(\debug_inst/vio0/vio_core_inst/word_count [11]), .I2(\debug_inst/vio0/vio_core_inst/word_count [10]), 
            .I3(\debug_inst/vio0/vio_core_inst/word_count [8]), .O(n4162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10324.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10325 (.I0(\debug_inst/vio0/vio_core_inst/word_count [15]), 
            .I1(\debug_inst/vio0/vio_core_inst/word_count [14]), .I2(\debug_inst/vio0/vio_core_inst/word_count [13]), 
            .I3(n4162), .O(n4163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10325.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10326 (.I0(\debug_inst/vio0/vio_core_inst/word_count [3]), 
            .I1(\debug_inst/vio0/vio_core_inst/word_count [2]), .I2(\debug_inst/vio0/vio_core_inst/word_count [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/word_count [0]), .O(n4164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10326.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10327 (.I0(n4163), .I1(n4159), .I2(n4164), .O(n4165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10327.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10328 (.I0(\debug_inst/vio0/vio_core_inst/word_count [15]), 
            .I1(\debug_inst/vio0/vio_core_inst/word_count [14]), .I2(\debug_inst/vio0/vio_core_inst/word_count [13]), 
            .I3(\debug_inst/vio0/vio_core_inst/word_count [9]), .O(n4166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10328.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10329 (.I0(n4158), .I1(n4159), .I2(n4162), .I3(n4166), 
            .O(n4167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10329.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10330 (.I0(n4167), .I1(n4150), .I2(n4137), .O(n4168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10330.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10331 (.I0(n4167), .I1(n4143), .I2(n4138), .I3(n4144), 
            .O(n4169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10331.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10332 (.I0(n4168), .I1(n4169), .I2(n4161), .I3(n4165), 
            .O(n4170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ee */ ;
    defparam LUT__10332.LUTMASK = 16'he0ee;
    EFX_LUT4 LUT__10333 (.I0(\debug_inst/vio0/vio_core_inst/module_state [1]), 
            .I1(\debug_inst/vio0/vio_core_inst/module_state [0]), .O(n4171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10333.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10334 (.I0(n4167), .I1(n4171), .I2(n4137), .O(n4172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10334.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10335 (.I0(n4144), .I1(n4149), .I2(n4143), .I3(n4153), 
            .O(n4173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__10335.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__10336 (.I0(n4170), .I1(n4152), .I2(n4172), .I3(n4173), 
            .O(\debug_inst/vio0/vio_core_inst/addr_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfeff */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1798)
    defparam LUT__10336.LUTMASK = 16'hfeff;
    EFX_LUT4 LUT__10337 (.I0(\debug_inst/edb_user_dr [45]), .I1(\debug_inst/vio0/vio_core_inst/word_count [0]), 
            .I2(n4139), .O(\debug_inst/vio0/vio_core_inst/data_to_word_counter [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1438)
    defparam LUT__10337.LUTMASK = 16'ha3a3;
    EFX_LUT4 LUT__10338 (.I0(n4123), .I1(bscan_CAPTURE), .I2(n4171), .O(n4174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__10338.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__10339 (.I0(n4155), .I1(\debug_inst/vio0/vio_core_inst/module_state [1]), 
            .I2(n4167), .I3(n4174), .O(n4175)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__10339.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__10340 (.I0(n4175), .I1(\debug_inst/vio0/vio_core_inst/module_state [0]), 
            .I2(n4144), .I3(n4154), .O(\debug_inst/vio0/vio_core_inst/word_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h10ff */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1798)
    defparam LUT__10340.LUTMASK = 16'h10ff;
    EFX_LUT4 LUT__10341 (.I0(\debug_inst/vio0/vio_core_inst/internal_register_select [0]), 
            .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [1]), 
            .I2(\debug_inst/vio0/vio_core_inst/internal_register_select [2]), 
            .O(n4176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9797 */ ;
    defparam LUT__10341.LUTMASK = 16'h9797;
    EFX_LUT4 LUT__10342 (.I0(n4123), .I1(bscan_CAPTURE), .O(n4177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10342.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10343 (.I0(n4139), .I1(n4177), .O(n4178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10343.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10344 (.I0(n4176), .I1(\debug_inst/vio0/vio_core_inst/data_from_biu [0]), 
            .I2(n4178), .O(n4179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__10344.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__10345 (.I0(\debug_inst/vio0/vio_core_inst/internal_register_select [0]), 
            .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [1]), 
            .I2(\debug_inst/vio0/vio_core_inst/internal_register_select [2]), 
            .O(n4180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10345.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10346 (.I0(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [0]), 
            .I1(n4180), .I2(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [1]), 
            .I3(n4178), .O(n4181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f */ ;
    defparam LUT__10346.LUTMASK = 16'h770f;
    EFX_LUT4 LUT__10347 (.I0(bscan_UPDATE), .I1(\debug_inst/vio0/vio_core_inst/module_state [1]), 
            .I2(\debug_inst/vio0/vio_core_inst/module_state [0]), .I3(\debug_inst/vio0/vio_core_inst/module_state [2]), 
            .O(n4182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__10347.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__10348 (.I0(\debug_inst/vio0/vio_core_inst/internal_register_select [3]), 
            .I1(n4182), .O(n4183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10348.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10349 (.I0(n4177), .I1(n4138), .I2(n4182), .I3(\debug_inst/vio0/vio_core_inst/module_state [3]), 
            .O(n4184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__10349.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__10350 (.I0(n4138), .I1(n4143), .I2(\debug_inst/vio0/vio_core_inst/module_state [2]), 
            .I3(n4184), .O(n4185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__10350.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__10351 (.I0(n4179), .I1(n4181), .I2(n4183), .I3(n4185), 
            .O(\debug_inst/vio0/vio_core_inst/n546 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a33 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam LUT__10351.LUTMASK = 16'h3a33;
    EFX_LUT4 LUT__10352 (.I0(\debug_inst/vio0/vio_core_inst/module_state [3]), 
            .I1(bscan_SHIFT), .I2(n4138), .O(n4186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10352.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10353 (.I0(\debug_inst/vio0/vio_core_inst/module_state [2]), 
            .I1(n4123), .I2(n4186), .I3(n4185), .O(ceg_net11)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__10353.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__10354 (.I0(\debug_inst/edb_user_dr [77]), .I1(\debug_inst/edb_user_dr [80]), 
            .I2(\debug_inst/edb_user_dr [78]), .I3(n4140), .O(\debug_inst/vio0/vio_core_inst/op_reg_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1798)
    defparam LUT__10354.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10355 (.I0(n4143), .I1(n4167), .I2(n4150), .O(n4187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__10355.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__10356 (.I0(bscan_UPDATE), .I1(n4167), .I2(n4138), .I3(n4143), 
            .O(n4188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10356.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10357 (.I0(n4188), .I1(n4187), .I2(n4175), .I3(n4144), 
            .O(n4189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10357.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10358 (.I0(\debug_inst/vio0/vio_core_inst/bit_count [4]), 
            .I1(\debug_inst/vio0/vio_core_inst/module_state [1]), .I2(\debug_inst/vio0/vio_core_inst/bit_count [5]), 
            .I3(n4115), .O(n4190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10358.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10359 (.I0(n4190), .I1(\debug_inst/vio0/vio_core_inst/module_state [0]), 
            .O(n4191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__10359.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__10360 (.I0(bscan_UPDATE), .I1(n4120), .O(n4192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10360.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10361 (.I0(\debug_inst/vio0/vio_core_inst/module_state [1]), 
            .I1(n4167), .I2(n4191), .I3(n4192), .O(n4193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__10361.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__10362 (.I0(n4177), .I1(n4114), .I2(n4137), .O(n4194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10362.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10363 (.I0(\debug_inst/vio0/vio_core_inst/op_reg_en ), .I1(n4189), 
            .I2(n4193), .I3(n4194), .O(\debug_inst/vio0/vio_core_inst/module_next_state [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfffe */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1613)
    defparam LUT__10363.LUTMASK = 16'hfffe;
    EFX_LUT4 LUT__10364 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [369]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [353]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10364.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10365 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [337]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [321]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4195), .O(n4196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10365.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10366 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [305]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [289]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10366.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10367 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [273]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [257]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4197), .O(n4198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10367.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10368 (.I0(n4198), .I1(n4196), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), .O(n4199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__10368.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__10369 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [113]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [97]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .O(n4200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__10369.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__10370 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [81]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [65]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .O(n4201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__10370.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__10371 (.I0(n4201), .I1(n4200), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), .O(n4202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__10371.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__10372 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [49]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [33]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .O(n4203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__10372.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__10373 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [17]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [1]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .O(n4204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__10373.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__10374 (.I0(n4204), .I1(n4203), .I2(\debug_inst/vio0/vio_core_inst/address_counter [3]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__10374.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__10375 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [241]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [225]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10375.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10376 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [209]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [193]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10376.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10377 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [177]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [161]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10377.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10378 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [145]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [129]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4208), .O(n4209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10378.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10379 (.I0(n4207), .I1(n4206), .I2(n4209), .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), 
            .O(n4210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__10379.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__10380 (.I0(n4205), .I1(n4202), .I2(n4210), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10380.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10381 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [497]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [481]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10381.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10382 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [465]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [449]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4212), .O(n4213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10382.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10383 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [433]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [417]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10383.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10384 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [401]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [385]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4214), .O(n4215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10384.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10385 (.I0(n4215), .I1(n4213), .I2(\debug_inst/vio0/vio_core_inst/address_counter [3]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), .O(n4216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__10385.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__10386 (.I0(n4199), .I1(n4216), .I2(n4211), .I3(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .O(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1836)
    defparam LUT__10386.LUTMASK = 16'h11f0;
    EFX_LUT4 LUT__10387 (.I0(\debug_inst/vio0/vio_core_inst/opcode [2]), .I1(\debug_inst/vio0/vio_core_inst/opcode [1]), 
            .O(n4217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10387.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10388 (.I0(n4170), .I1(n4172), .I2(n4173), .I3(n4217), 
            .O(\debug_inst/vio0/vio_core_inst/n2907 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1839)
    defparam LUT__10388.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10389 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [368]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [352]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10389.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10390 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [336]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [320]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4218), .O(n4219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10390.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10391 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [304]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [288]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10391.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10392 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [272]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [256]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4220), .O(n4221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10392.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10393 (.I0(n4221), .I1(n4219), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), .O(n4222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__10393.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__10394 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [112]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [96]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .O(n4223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__10394.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__10395 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [80]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [64]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .O(n4224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__10395.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__10396 (.I0(n4224), .I1(n4223), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), .O(n4225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__10396.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__10397 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [48]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [32]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .O(n4226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__10397.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__10398 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [16]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [0]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .O(n4227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__10398.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__10399 (.I0(n4227), .I1(n4226), .I2(\debug_inst/vio0/vio_core_inst/address_counter [3]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__10399.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__10400 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [240]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [224]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10400.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10401 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [208]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [192]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10401.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10402 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [176]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [160]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10402.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10403 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [144]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [128]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4231), .O(n4232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10403.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10404 (.I0(n4230), .I1(n4229), .I2(n4232), .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), 
            .O(n4233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f */ ;
    defparam LUT__10404.LUTMASK = 16'hee0f;
    EFX_LUT4 LUT__10405 (.I0(n4228), .I1(n4225), .I2(n4233), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10405.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10406 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [496]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [480]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10406.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10407 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [464]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [448]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4235), .O(n4236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10407.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10408 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [432]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [416]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10408.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10409 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [400]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [384]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4237), .O(n4238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10409.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10410 (.I0(n4238), .I1(n4236), .I2(\debug_inst/vio0/vio_core_inst/address_counter [3]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), .O(n4239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__10410.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__10411 (.I0(n4222), .I1(n4239), .I2(n4234), .I3(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .O(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1836)
    defparam LUT__10411.LUTMASK = 16'h11f0;
    EFX_LUT4 LUT__10412 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [383]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [367]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10412.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10413 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [351]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [335]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10413.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10414 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [511]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [495]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10414.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10415 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [479]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [463]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10415.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10416 (.I0(n4242), .I1(n4243), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10416.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10417 (.I0(n4241), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4240), .I3(n4244), .O(n4245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10417.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10418 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [319]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [303]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10418.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10419 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [287]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [271]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10419.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10420 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [447]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [431]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10420.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10421 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [415]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [399]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10421.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10422 (.I0(n4248), .I1(n4249), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10422.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10423 (.I0(n4247), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4246), .I3(n4250), .O(n4251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10423.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10424 (.I0(n4245), .I1(n4251), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), .O(n4252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10424.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10425 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [255]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [239]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10425.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10426 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [223]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [207]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10426.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10427 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [127]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [111]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10427.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10428 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [95]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [79]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4255), .O(n4256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10428.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10429 (.I0(n4254), .I1(n4253), .I2(n4256), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10429.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10430 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [31]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [15]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10430.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10431 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [63]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [47]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10431.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10432 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [191]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [175]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10432.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10433 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [159]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [143]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4260), .O(n4261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10433.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10434 (.I0(n4259), .I1(n4258), .I2(n4261), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10434.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10435 (.I0(n4262), .I1(n4257), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(n4252), .O(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1836)
    defparam LUT__10435.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__10436 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [382]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [366]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10436.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10437 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [350]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [334]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10437.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10438 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [510]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [494]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10438.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10439 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [478]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [462]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10439.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10440 (.I0(n4265), .I1(n4266), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10440.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10441 (.I0(n4264), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4263), .I3(n4267), .O(n4268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10441.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10442 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [318]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [302]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10442.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10443 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [286]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [270]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10443.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10444 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [446]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [430]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10444.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10445 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [414]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [398]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10445.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10446 (.I0(n4271), .I1(n4272), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10446.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10447 (.I0(n4270), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4269), .I3(n4273), .O(n4274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10447.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10448 (.I0(n4268), .I1(n4274), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), .O(n4275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10448.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10449 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [254]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [238]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10449.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10450 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [222]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [206]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10450.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10451 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [126]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [110]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10451.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10452 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [94]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [78]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4278), .O(n4279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10452.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10453 (.I0(n4277), .I1(n4276), .I2(n4279), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10453.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10454 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [30]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [14]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10454.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10455 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [62]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [46]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10455.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10456 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [190]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [174]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10456.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10457 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [158]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [142]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4283), .O(n4284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10457.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10458 (.I0(n4282), .I1(n4281), .I2(n4284), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10458.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10459 (.I0(n4285), .I1(n4280), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(n4275), .O(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1836)
    defparam LUT__10459.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__10460 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [381]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [365]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10460.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10461 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [349]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [333]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10461.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10462 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [509]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [493]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10462.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10463 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [477]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [461]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10463.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10464 (.I0(n4288), .I1(n4289), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10464.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10465 (.I0(n4287), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4286), .I3(n4290), .O(n4291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10465.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10466 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [317]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [301]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10466.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10467 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [285]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [269]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10467.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10468 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [445]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [429]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10468.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10469 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [413]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [397]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10469.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10470 (.I0(n4294), .I1(n4295), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10470.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10471 (.I0(n4293), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4292), .I3(n4296), .O(n4297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10471.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10472 (.I0(n4291), .I1(n4297), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), .O(n4298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10472.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10473 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [253]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [237]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10473.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10474 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [221]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [205]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10474.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10475 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [125]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [109]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10475.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10476 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [93]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [77]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4301), .O(n4302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10476.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10477 (.I0(n4300), .I1(n4299), .I2(n4302), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10477.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10478 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [29]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [13]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10478.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10479 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [61]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [45]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10479.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10480 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [189]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [173]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10480.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10481 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [157]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [141]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4306), .O(n4307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10481.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10482 (.I0(n4305), .I1(n4304), .I2(n4307), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10482.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10483 (.I0(n4308), .I1(n4303), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(n4298), .O(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1836)
    defparam LUT__10483.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__10484 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [380]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [364]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10484.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10485 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [348]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [332]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10485.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10486 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [508]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [492]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10486.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10487 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [476]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [460]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10487.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10488 (.I0(n4311), .I1(n4312), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10488.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10489 (.I0(n4310), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4309), .I3(n4313), .O(n4314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10489.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10490 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [316]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [300]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10490.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10491 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [284]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [268]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10491.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10492 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [444]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [428]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10492.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10493 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [412]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [396]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10493.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10494 (.I0(n4317), .I1(n4318), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10494.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10495 (.I0(n4316), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4315), .I3(n4319), .O(n4320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10495.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10496 (.I0(n4314), .I1(n4320), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), .O(n4321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10496.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10497 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [252]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [236]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10497.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10498 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [220]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [204]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10498.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10499 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [124]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [108]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10499.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10500 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [92]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [76]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4324), .O(n4325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10500.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10501 (.I0(n4323), .I1(n4322), .I2(n4325), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10501.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10502 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [28]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [12]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10502.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10503 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [60]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [44]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10503.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10504 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [188]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [172]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10504.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10505 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [156]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [140]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4329), .O(n4330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10505.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10506 (.I0(n4328), .I1(n4327), .I2(n4330), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10506.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10507 (.I0(n4331), .I1(n4326), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(n4321), .O(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1836)
    defparam LUT__10507.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__10508 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [379]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [363]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10508.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10509 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [347]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [331]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10509.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10510 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [507]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [491]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10510.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10511 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [475]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [459]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10511.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10512 (.I0(n4334), .I1(n4335), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10512.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10513 (.I0(n4333), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4332), .I3(n4336), .O(n4337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10513.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10514 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [315]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [299]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10514.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10515 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [283]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [267]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10515.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10516 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [443]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [427]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10516.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10517 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [411]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [395]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10517.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10518 (.I0(n4340), .I1(n4341), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10518.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10519 (.I0(n4339), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4338), .I3(n4342), .O(n4343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10519.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10520 (.I0(n4337), .I1(n4343), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), .O(n4344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10520.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10521 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [251]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [235]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10521.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10522 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [219]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [203]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10522.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10523 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [123]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [107]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10523.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10524 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [91]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [75]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4347), .O(n4348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10524.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10525 (.I0(n4346), .I1(n4345), .I2(n4348), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10525.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10526 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [27]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [11]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10526.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10527 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [59]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [43]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10527.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10528 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [187]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [171]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10528.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10529 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [155]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [139]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4352), .O(n4353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10529.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10530 (.I0(n4351), .I1(n4350), .I2(n4353), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10530.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10531 (.I0(n4354), .I1(n4349), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(n4344), .O(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1836)
    defparam LUT__10531.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__10532 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [378]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [362]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10532.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10533 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [346]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [330]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10533.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10534 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [506]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [490]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10534.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10535 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [474]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [458]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10535.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10536 (.I0(n4357), .I1(n4358), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10536.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10537 (.I0(n4356), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4355), .I3(n4359), .O(n4360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10537.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10538 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [314]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [298]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10538.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10539 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [282]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [266]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10539.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10540 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [442]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [426]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10540.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10541 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [410]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [394]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10541.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10542 (.I0(n4363), .I1(n4364), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10542.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10543 (.I0(n4362), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4361), .I3(n4365), .O(n4366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10543.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10544 (.I0(n4360), .I1(n4366), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), .O(n4367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10544.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10545 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [250]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [234]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10545.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10546 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [218]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [202]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10546.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10547 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [122]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [106]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10547.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10548 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [90]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [74]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4370), .O(n4371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10548.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10549 (.I0(n4369), .I1(n4368), .I2(n4371), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10549.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10550 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [26]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [10]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10550.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10551 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [58]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [42]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10551.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10552 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [186]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [170]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10552.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10553 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [154]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [138]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4375), .O(n4376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10553.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10554 (.I0(n4374), .I1(n4373), .I2(n4376), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10554.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10555 (.I0(n4377), .I1(n4372), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(n4367), .O(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1836)
    defparam LUT__10555.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__10556 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [377]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [361]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10556.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10557 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [345]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [329]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10557.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10558 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [505]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [489]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10558.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10559 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [473]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [457]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10559.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10560 (.I0(n4380), .I1(n4381), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10560.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10561 (.I0(n4379), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4378), .I3(n4382), .O(n4383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10561.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10562 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [313]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [297]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10562.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10563 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [281]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [265]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10563.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10564 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [441]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [425]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10564.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10565 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [409]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [393]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10565.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10566 (.I0(n4386), .I1(n4387), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10566.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10567 (.I0(n4385), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4384), .I3(n4388), .O(n4389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10567.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10568 (.I0(n4383), .I1(n4389), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), .O(n4390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10568.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10569 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [249]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [233]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10569.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10570 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [217]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [201]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10570.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10571 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [121]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [105]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10571.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10572 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [89]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [73]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4393), .O(n4394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10572.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10573 (.I0(n4392), .I1(n4391), .I2(n4394), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10573.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10574 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [25]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [9]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10574.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10575 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [57]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [41]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10575.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10576 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [185]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [169]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10576.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10577 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [153]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [137]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4398), .O(n4399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10577.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10578 (.I0(n4397), .I1(n4396), .I2(n4399), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10578.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10579 (.I0(n4400), .I1(n4395), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(n4390), .O(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1836)
    defparam LUT__10579.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__10580 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [376]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [360]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10580.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10581 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [344]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [328]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10581.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10582 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [504]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [488]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10582.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10583 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [472]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [456]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10583.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10584 (.I0(n4403), .I1(n4404), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10584.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10585 (.I0(n4402), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4401), .I3(n4405), .O(n4406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10585.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10586 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [312]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [296]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10586.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10587 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [280]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [264]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10587.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10588 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [440]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [424]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10588.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10589 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [408]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [392]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10589.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10590 (.I0(n4409), .I1(n4410), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10590.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10591 (.I0(n4408), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4407), .I3(n4411), .O(n4412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10591.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10592 (.I0(n4406), .I1(n4412), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), .O(n4413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10592.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10593 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [248]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [232]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10593.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10594 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [216]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [200]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10594.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10595 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [120]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [104]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10595.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10596 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [88]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [72]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4416), .O(n4417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10596.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10597 (.I0(n4415), .I1(n4414), .I2(n4417), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10597.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10598 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [24]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [8]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10598.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10599 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [56]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [40]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10599.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10600 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [184]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [168]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10600.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10601 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [152]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [136]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4421), .O(n4422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10601.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10602 (.I0(n4420), .I1(n4419), .I2(n4422), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10602.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10603 (.I0(n4423), .I1(n4418), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(n4413), .O(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1836)
    defparam LUT__10603.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__10604 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [375]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [359]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10604.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10605 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [343]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [327]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10605.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10606 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [503]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [487]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10606.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10607 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [471]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [455]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10607.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10608 (.I0(n4426), .I1(n4427), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10608.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10609 (.I0(n4425), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4424), .I3(n4428), .O(n4429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10609.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10610 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [311]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [295]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10610.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10611 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [279]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [263]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10611.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10612 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [439]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [423]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10612.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10613 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [407]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [391]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10613.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10614 (.I0(n4432), .I1(n4433), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10614.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10615 (.I0(n4431), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4430), .I3(n4434), .O(n4435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10615.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10616 (.I0(n4429), .I1(n4435), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), .O(n4436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10616.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10617 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [247]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [231]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10617.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10618 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [215]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [199]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10618.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10619 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [119]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [103]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10619.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10620 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [87]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [71]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4439), .O(n4440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10620.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10621 (.I0(n4438), .I1(n4437), .I2(n4440), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10621.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10622 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [23]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [7]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10622.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10623 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [55]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [39]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10623.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10624 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [183]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [167]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10624.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10625 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [151]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [135]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4444), .O(n4445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10625.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10626 (.I0(n4443), .I1(n4442), .I2(n4445), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10626.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10627 (.I0(n4446), .I1(n4441), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(n4436), .O(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1836)
    defparam LUT__10627.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__10628 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [374]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [358]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10628.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10629 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [342]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [326]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10629.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10630 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [502]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [486]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10630.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10631 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [470]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [454]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10631.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10632 (.I0(n4449), .I1(n4450), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10632.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10633 (.I0(n4448), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4447), .I3(n4451), .O(n4452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10633.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10634 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [310]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [294]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10634.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10635 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [278]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [262]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10635.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10636 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [438]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [422]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10636.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10637 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [406]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [390]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10637.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10638 (.I0(n4455), .I1(n4456), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10638.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10639 (.I0(n4454), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4453), .I3(n4457), .O(n4458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10639.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10640 (.I0(n4452), .I1(n4458), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), .O(n4459)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10640.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10641 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [246]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [230]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10641.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10642 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [214]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [198]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10642.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10643 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [118]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [102]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10643.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10644 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [86]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [70]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4462), .O(n4463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10644.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10645 (.I0(n4461), .I1(n4460), .I2(n4463), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10645.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10646 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [22]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [6]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10646.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10647 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [54]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [38]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10647.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10648 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [182]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [166]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10648.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10649 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [150]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [134]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4467), .O(n4468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10649.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10650 (.I0(n4466), .I1(n4465), .I2(n4468), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10650.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10651 (.I0(n4469), .I1(n4464), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(n4459), .O(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1836)
    defparam LUT__10651.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__10652 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [373]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [357]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10652.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10653 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [341]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [325]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10653.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10654 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [501]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [485]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10654.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10655 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [469]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [453]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10655.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10656 (.I0(n4472), .I1(n4473), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10656.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10657 (.I0(n4471), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4470), .I3(n4474), .O(n4475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10657.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10658 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [309]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [293]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10658.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10659 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [277]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [261]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10659.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10660 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [437]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [421]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10660.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10661 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [405]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [389]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10661.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10662 (.I0(n4478), .I1(n4479), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10662.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10663 (.I0(n4477), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4476), .I3(n4480), .O(n4481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10663.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10664 (.I0(n4475), .I1(n4481), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), .O(n4482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10664.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10665 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [245]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [229]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10665.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10666 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [213]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [197]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10666.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10667 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [117]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [101]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10667.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10668 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [85]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [69]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4485), .O(n4486)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10668.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10669 (.I0(n4484), .I1(n4483), .I2(n4486), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10669.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10670 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [21]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [5]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10670.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10671 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [53]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [37]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10671.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10672 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [181]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [165]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10672.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10673 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [149]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [133]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4490), .O(n4491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10673.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10674 (.I0(n4489), .I1(n4488), .I2(n4491), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4492)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10674.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10675 (.I0(n4492), .I1(n4487), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(n4482), .O(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1836)
    defparam LUT__10675.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__10676 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [372]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [356]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10676.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10677 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [340]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [324]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10677.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10678 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [500]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [484]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10678.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10679 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [468]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [452]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10679.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10680 (.I0(n4495), .I1(n4496), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10680.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10681 (.I0(n4494), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4493), .I3(n4497), .O(n4498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10681.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10682 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [308]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [292]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10682.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10683 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [276]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [260]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10683.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10684 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [436]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [420]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10684.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10685 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [404]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [388]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10685.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10686 (.I0(n4501), .I1(n4502), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10686.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10687 (.I0(n4500), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4499), .I3(n4503), .O(n4504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10687.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10688 (.I0(n4498), .I1(n4504), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), .O(n4505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10688.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10689 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [244]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [228]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10689.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10690 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [212]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [196]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10690.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10691 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [116]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [100]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10691.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10692 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [84]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [68]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4508), .O(n4509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10692.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10693 (.I0(n4507), .I1(n4506), .I2(n4509), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10693.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10694 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [20]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [4]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10694.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10695 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [52]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [36]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10695.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10696 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [180]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [164]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10696.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10697 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [148]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [132]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4513), .O(n4514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10697.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10698 (.I0(n4512), .I1(n4511), .I2(n4514), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10698.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10699 (.I0(n4515), .I1(n4510), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(n4505), .O(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1836)
    defparam LUT__10699.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__10700 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [371]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [355]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10700.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10701 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [339]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [323]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10701.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10702 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [499]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [483]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10702.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10703 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [467]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [451]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10703.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10704 (.I0(n4518), .I1(n4519), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10704.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10705 (.I0(n4517), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4516), .I3(n4520), .O(n4521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10705.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10706 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [307]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [291]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4522)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10706.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10707 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [275]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [259]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10707.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10708 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [435]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [419]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10708.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10709 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [403]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [387]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10709.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10710 (.I0(n4524), .I1(n4525), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10710.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10711 (.I0(n4523), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4522), .I3(n4526), .O(n4527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10711.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10712 (.I0(n4521), .I1(n4527), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), .O(n4528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10712.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10713 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [243]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [227]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10713.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10714 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [211]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [195]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10714.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10715 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [115]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [99]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10715.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10716 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [83]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [67]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4531), .O(n4532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10716.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10717 (.I0(n4530), .I1(n4529), .I2(n4532), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10717.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10718 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [19]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [3]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10718.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10719 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [51]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [35]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10719.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10720 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [179]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [163]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10720.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10721 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [147]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [131]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4536), .O(n4537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10721.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10722 (.I0(n4535), .I1(n4534), .I2(n4537), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10722.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10723 (.I0(n4538), .I1(n4533), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(n4528), .O(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1836)
    defparam LUT__10723.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__10724 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [370]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [354]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10724.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10725 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [338]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [322]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10725.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10726 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [498]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [482]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10726.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10727 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [466]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [450]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10727.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10728 (.I0(n4541), .I1(n4542), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10728.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10729 (.I0(n4540), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4539), .I3(n4543), .O(n4544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10729.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10730 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [306]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [290]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10730.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10731 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [274]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [258]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10731.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10732 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [434]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [418]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__10732.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__10733 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [402]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [386]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__10733.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__10734 (.I0(n4547), .I1(n4548), .I2(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10734.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10735 (.I0(n4546), .I1(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .I2(n4545), .I3(n4549), .O(n4550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe */ ;
    defparam LUT__10735.LUTMASK = 16'h00fe;
    EFX_LUT4 LUT__10736 (.I0(n4544), .I1(n4550), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [3]), .O(n4551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10736.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10737 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [242]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [226]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10737.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10738 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [210]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [194]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10738.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10739 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [114]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [98]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10739.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10740 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [82]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [66]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4554), .O(n4555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__10740.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__10741 (.I0(n4553), .I1(n4552), .I2(n4555), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10741.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10742 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [18]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [2]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__10742.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__10743 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [50]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [34]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [2]), .O(n4558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10743.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10744 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [178]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [162]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/address_counter [1]), .O(n4559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10744.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10745 (.I0(\debug_inst/vio0/vio_core_inst/probe_in_sync [146]), 
            .I1(\debug_inst/vio0/vio_core_inst/probe_in_sync [130]), .I2(\debug_inst/vio0/vio_core_inst/address_counter [2]), 
            .I3(n4559), .O(n4560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10745.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10746 (.I0(n4558), .I1(n4557), .I2(n4560), .I3(\debug_inst/vio0/vio_core_inst/address_counter [4]), 
            .O(n4561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10746.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10747 (.I0(n4561), .I1(n4556), .I2(\debug_inst/vio0/vio_core_inst/address_counter [5]), 
            .I3(n4551), .O(\debug_inst/vio0/vio_core_inst/probe_in_mux_out [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1836)
    defparam LUT__10747.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__10748 (.I0(bscan_TDI), .I1(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [0]), 
            .I2(\debug_inst/vio0/vio_core_inst/module_state [1]), .I3(\debug_inst/vio0/vio_core_inst/crc_data_out [0]), 
            .O(n4562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h53ac */ ;
    defparam LUT__10748.LUTMASK = 16'h53ac;
    EFX_LUT4 LUT__10749 (.I0(n4562), .I1(n4156), .O(n4563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10749.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10750 (.I0(n4563), .I1(n4152), .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10750.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10751 (.I0(n4171), .I1(n4120), .O(n4564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10751.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10752 (.I0(n4564), .I1(bscan_SHIFT), .I2(n4152), .I3(n4156), 
            .O(ceg_net16)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(307)
    defparam LUT__10752.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__10753 (.I0(n4152), .I1(n4563), .I2(\debug_inst/vio0/vio_core_inst/crc_data_out [31]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10753.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__10754 (.I0(n4152), .I1(n4563), .I2(\debug_inst/vio0/vio_core_inst/crc_data_out [30]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10754.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__10755 (.I0(n4152), .I1(\debug_inst/vio0/vio_core_inst/crc_data_out [29]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10755.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10756 (.I0(n4152), .I1(n4563), .I2(\debug_inst/vio0/vio_core_inst/crc_data_out [28]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10756.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__10757 (.I0(n4152), .I1(n4563), .I2(\debug_inst/vio0/vio_core_inst/crc_data_out [27]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10757.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__10758 (.I0(n4152), .I1(\debug_inst/vio0/vio_core_inst/crc_data_out [26]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10758.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10759 (.I0(n4152), .I1(n4563), .I2(\debug_inst/vio0/vio_core_inst/crc_data_out [25]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10759.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__10760 (.I0(n4152), .I1(n4563), .I2(\debug_inst/vio0/vio_core_inst/crc_data_out [24]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10760.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__10761 (.I0(n4152), .I1(\debug_inst/vio0/vio_core_inst/crc_data_out [23]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10761.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10762 (.I0(n4152), .I1(n4563), .I2(\debug_inst/vio0/vio_core_inst/crc_data_out [22]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10762.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__10763 (.I0(n4152), .I1(n4563), .I2(\debug_inst/vio0/vio_core_inst/crc_data_out [21]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10763.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__10764 (.I0(n4152), .I1(n4563), .I2(\debug_inst/vio0/vio_core_inst/crc_data_out [20]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10764.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__10765 (.I0(n4152), .I1(\debug_inst/vio0/vio_core_inst/crc_data_out [19]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10765.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10766 (.I0(n4152), .I1(\debug_inst/vio0/vio_core_inst/crc_data_out [18]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10766.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10767 (.I0(n4152), .I1(\debug_inst/vio0/vio_core_inst/crc_data_out [17]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10767.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10768 (.I0(n4152), .I1(n4563), .I2(\debug_inst/vio0/vio_core_inst/crc_data_out [16]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10768.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__10769 (.I0(n4152), .I1(\debug_inst/vio0/vio_core_inst/crc_data_out [15]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10769.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10770 (.I0(n4152), .I1(\debug_inst/vio0/vio_core_inst/crc_data_out [14]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10770.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10771 (.I0(n4152), .I1(\debug_inst/vio0/vio_core_inst/crc_data_out [13]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10771.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10772 (.I0(n4152), .I1(\debug_inst/vio0/vio_core_inst/crc_data_out [12]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10772.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10773 (.I0(n4152), .I1(\debug_inst/vio0/vio_core_inst/crc_data_out [11]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10773.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10774 (.I0(n4152), .I1(n4563), .I2(\debug_inst/vio0/vio_core_inst/crc_data_out [10]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10774.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__10775 (.I0(n4152), .I1(n4563), .I2(\debug_inst/vio0/vio_core_inst/crc_data_out [9]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10775.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__10776 (.I0(n4152), .I1(\debug_inst/vio0/vio_core_inst/crc_data_out [8]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10776.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10777 (.I0(n4152), .I1(\debug_inst/vio0/vio_core_inst/crc_data_out [7]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10777.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10778 (.I0(n4152), .I1(n4563), .I2(\debug_inst/vio0/vio_core_inst/crc_data_out [6]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10778.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__10779 (.I0(n4152), .I1(\debug_inst/vio0/vio_core_inst/crc_data_out [5]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10779.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10780 (.I0(n4152), .I1(\debug_inst/vio0/vio_core_inst/crc_data_out [4]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10780.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10781 (.I0(n4152), .I1(\debug_inst/vio0/vio_core_inst/crc_data_out [3]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10781.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10782 (.I0(n4152), .I1(\debug_inst/vio0/vio_core_inst/crc_data_out [2]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10782.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10783 (.I0(n4152), .I1(\debug_inst/vio0/vio_core_inst/crc_data_out [1]), 
            .O(\debug_inst/vio0/vio_core_inst/axi_crc_i/n118 [0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(361)
    defparam LUT__10783.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10784 (.I0(n4167), .I1(n4138), .I2(n4192), .O(n4565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__10784.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__10785 (.I0(bscan_UPDATE), .I1(n4145), .I2(n4167), .I3(n4565), 
            .O(\debug_inst/vio0/vio_core_inst/module_next_state [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1613)
    defparam LUT__10785.LUTMASK = 16'hff40;
    EFX_LUT4 LUT__10786 (.I0(n4143), .I1(\debug_inst/vio0/vio_core_inst/module_state [0]), 
            .I2(\debug_inst/vio0/vio_core_inst/module_state [1]), .I3(n4144), 
            .O(n4566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7100 */ ;
    defparam LUT__10786.LUTMASK = 16'h7100;
    EFX_LUT4 LUT__10787 (.I0(n4153), .I1(n4171), .I2(bscan_UPDATE), .I3(n4144), 
            .O(n4567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcf0a */ ;
    defparam LUT__10787.LUTMASK = 16'hcf0a;
    EFX_LUT4 LUT__10788 (.I0(n4566), .I1(n4167), .I2(n4567), .I3(n4151), 
            .O(\debug_inst/vio0/vio_core_inst/module_next_state [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffb0 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1613)
    defparam LUT__10788.LUTMASK = 16'hffb0;
    EFX_LUT4 LUT__10789 (.I0(bscan_UPDATE), .I1(\debug_inst/vio0/vio_core_inst/module_state [0]), 
            .I2(\debug_inst/vio0/vio_core_inst/module_state [2]), .I3(\debug_inst/vio0/vio_core_inst/module_state [1]), 
            .O(n4568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__10789.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__10790 (.I0(n4177), .I1(\debug_inst/vio0/vio_core_inst/module_state [2]), 
            .I2(n4167), .I3(n4171), .O(n4569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__10790.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__10791 (.I0(n4569), .I1(n4568), .I2(\debug_inst/vio0/vio_core_inst/module_state [3]), 
            .O(n4570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__10791.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__10792 (.I0(n4171), .I1(n4192), .I2(n4570), .O(\debug_inst/vio0/vio_core_inst/module_next_state [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1613)
    defparam LUT__10792.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__10793 (.I0(\debug_inst/vio0/vio_core_inst/internal_register_select [3]), 
            .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [1]), 
            .I2(\debug_inst/vio0/vio_core_inst/data_from_biu [15]), .I3(n4182), 
            .O(n4571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f */ ;
    defparam LUT__10793.LUTMASK = 16'h770f;
    EFX_LUT4 LUT__10794 (.I0(n4571), .I1(n4185), .O(\debug_inst/vio0/vio_core_inst/n546 [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam LUT__10794.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10795 (.I0(\debug_inst/vio0/vio_core_inst/internal_register_select [0]), 
            .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [2]), 
            .I2(\debug_inst/vio0/vio_core_inst/internal_register_select [1]), 
            .O(n4572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__10795.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__10796 (.I0(n4572), .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [3]), 
            .I2(\debug_inst/vio0/vio_core_inst/data_from_biu [14]), .I3(n4182), 
            .O(n4573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__10796.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__10797 (.I0(n4573), .I1(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [15]), 
            .I2(n4185), .O(\debug_inst/vio0/vio_core_inst/n546 [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam LUT__10797.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__10798 (.I0(\debug_inst/vio0/vio_core_inst/internal_register_select [0]), 
            .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [1]), 
            .I2(\debug_inst/vio0/vio_core_inst/internal_register_select [2]), 
            .O(n4574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__10798.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__10799 (.I0(n4574), .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [3]), 
            .I2(\debug_inst/vio0/vio_core_inst/data_from_biu [13]), .I3(n4182), 
            .O(n4575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__10799.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__10800 (.I0(n4575), .I1(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [14]), 
            .I2(n4185), .O(\debug_inst/vio0/vio_core_inst/n546 [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam LUT__10800.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__10801 (.I0(\debug_inst/vio0/vio_core_inst/internal_register_select [1]), 
            .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [2]), 
            .I2(\debug_inst/vio0/vio_core_inst/internal_register_select [0]), 
            .I3(\debug_inst/vio0/vio_core_inst/internal_register_select [3]), 
            .O(n4576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__10801.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__10802 (.I0(\debug_inst/vio0/vio_core_inst/internal_register_select [1]), 
            .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [2]), 
            .I2(n4576), .O(n4577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__10802.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__10803 (.I0(n4577), .I1(\debug_inst/vio0/vio_core_inst/data_from_biu [12]), 
            .I2(n4182), .O(n4578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__10803.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__10804 (.I0(n4578), .I1(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [13]), 
            .I2(n4185), .O(\debug_inst/vio0/vio_core_inst/n546 [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam LUT__10804.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__10805 (.I0(\debug_inst/vio0/vio_core_inst/internal_register_select [0]), 
            .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [2]), 
            .I2(\debug_inst/vio0/vio_core_inst/internal_register_select [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/internal_register_select [3]), 
            .O(n4579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__10805.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__10806 (.I0(n4579), .I1(\debug_inst/vio0/vio_core_inst/data_from_biu [11]), 
            .I2(n4182), .O(n4580)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__10806.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__10807 (.I0(n4580), .I1(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [12]), 
            .I2(n4185), .O(\debug_inst/vio0/vio_core_inst/n546 [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam LUT__10807.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__10808 (.I0(\debug_inst/vio0/vio_core_inst/internal_register_select [0]), 
            .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [2]), 
            .I2(\debug_inst/vio0/vio_core_inst/internal_register_select [1]), 
            .O(n4581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;
    defparam LUT__10808.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__10809 (.I0(n4581), .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [3]), 
            .I2(\debug_inst/vio0/vio_core_inst/data_from_biu [10]), .I3(n4182), 
            .O(n4582)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__10809.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__10810 (.I0(n4582), .I1(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [11]), 
            .I2(n4185), .O(\debug_inst/vio0/vio_core_inst/n546 [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam LUT__10810.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__10811 (.I0(n4576), .I1(\debug_inst/vio0/vio_core_inst/data_from_biu [9]), 
            .I2(n4182), .O(n4583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__10811.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__10812 (.I0(n4583), .I1(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [10]), 
            .I2(n4185), .O(\debug_inst/vio0/vio_core_inst/n546 [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam LUT__10812.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__10813 (.I0(\debug_inst/vio0/vio_core_inst/internal_register_select [0]), 
            .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [1]), 
            .I2(\debug_inst/vio0/vio_core_inst/internal_register_select [2]), 
            .I3(\debug_inst/vio0/vio_core_inst/internal_register_select [3]), 
            .O(n4584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4200 */ ;
    defparam LUT__10813.LUTMASK = 16'h4200;
    EFX_LUT4 LUT__10814 (.I0(n4584), .I1(\debug_inst/vio0/vio_core_inst/data_from_biu [8]), 
            .I2(n4182), .O(n4585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__10814.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__10815 (.I0(n4585), .I1(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [9]), 
            .I2(n4185), .O(\debug_inst/vio0/vio_core_inst/n546 [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam LUT__10815.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__10816 (.I0(\debug_inst/vio0/vio_core_inst/internal_register_select [2]), 
            .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [1]), 
            .I2(\debug_inst/vio0/vio_core_inst/internal_register_select [0]), 
            .O(n4586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;
    defparam LUT__10816.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__10817 (.I0(n4586), .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [3]), 
            .I2(\debug_inst/vio0/vio_core_inst/data_from_biu [7]), .I3(n4182), 
            .O(n4587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__10817.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__10818 (.I0(n4587), .I1(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [8]), 
            .I2(n4185), .O(\debug_inst/vio0/vio_core_inst/n546 [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam LUT__10818.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__10819 (.I0(\debug_inst/vio0/vio_core_inst/internal_register_select [1]), 
            .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [0]), 
            .I2(\debug_inst/vio0/vio_core_inst/internal_register_select [2]), 
            .O(n4588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b */ ;
    defparam LUT__10819.LUTMASK = 16'h4b4b;
    EFX_LUT4 LUT__10820 (.I0(\debug_inst/vio0/vio_core_inst/internal_register_select [3]), 
            .I1(n4588), .I2(\debug_inst/vio0/vio_core_inst/data_from_biu [6]), 
            .I3(n4182), .O(n4589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f */ ;
    defparam LUT__10820.LUTMASK = 16'h770f;
    EFX_LUT4 LUT__10821 (.I0(n4589), .I1(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [7]), 
            .I2(n4185), .O(\debug_inst/vio0/vio_core_inst/n546 [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam LUT__10821.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__10822 (.I0(\debug_inst/vio0/vio_core_inst/internal_register_select [3]), 
            .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [2]), 
            .I2(\debug_inst/vio0/vio_core_inst/internal_register_select [0]), 
            .I3(\debug_inst/vio0/vio_core_inst/internal_register_select [1]), 
            .O(n4590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha82a */ ;
    defparam LUT__10822.LUTMASK = 16'ha82a;
    EFX_LUT4 LUT__10823 (.I0(n4590), .I1(\debug_inst/vio0/vio_core_inst/data_from_biu [5]), 
            .I2(n4182), .O(n4591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__10823.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__10824 (.I0(n4591), .I1(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [6]), 
            .I2(n4185), .O(\debug_inst/vio0/vio_core_inst/n546 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam LUT__10824.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__10825 (.I0(\debug_inst/vio0/vio_core_inst/internal_register_select [2]), 
            .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [1]), 
            .I2(\debug_inst/vio0/vio_core_inst/internal_register_select [0]), 
            .O(n4592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;
    defparam LUT__10825.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__10826 (.I0(n4592), .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [3]), 
            .I2(\debug_inst/vio0/vio_core_inst/data_from_biu [4]), .I3(n4182), 
            .O(n4593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__10826.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__10827 (.I0(n4593), .I1(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [5]), 
            .I2(n4185), .O(\debug_inst/vio0/vio_core_inst/n546 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam LUT__10827.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__10828 (.I0(n4574), .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [3]), 
            .I2(\debug_inst/vio0/vio_core_inst/data_from_biu [3]), .I3(n4182), 
            .O(n4594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__10828.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__10829 (.I0(n4594), .I1(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [4]), 
            .I2(n4185), .O(\debug_inst/vio0/vio_core_inst/n546 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam LUT__10829.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__10830 (.I0(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [2]), 
            .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [1]), 
            .I2(\debug_inst/vio0/vio_core_inst/internal_register_select [2]), 
            .I3(n4183), .O(n4595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfdc3 */ ;
    defparam LUT__10830.LUTMASK = 16'hfdc3;
    EFX_LUT4 LUT__10831 (.I0(\debug_inst/vio0/vio_core_inst/internal_register_select [0]), 
            .I1(n4595), .I2(\debug_inst/vio0/vio_core_inst/data_from_biu [2]), 
            .I3(n4178), .O(n4596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10831.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10832 (.I0(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [3]), 
            .I1(n4178), .I2(n4596), .I3(n4185), .O(\debug_inst/vio0/vio_core_inst/n546 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3cae */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam LUT__10832.LUTMASK = 16'h3cae;
    EFX_LUT4 LUT__10833 (.I0(\debug_inst/vio0/vio_core_inst/internal_register_select [0]), 
            .I1(\debug_inst/vio0/vio_core_inst/internal_register_select [1]), 
            .I2(\debug_inst/vio0/vio_core_inst/internal_register_select [2]), 
            .O(n4597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__10833.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__10834 (.I0(\debug_inst/vio0/vio_core_inst/internal_reg_r0 [1]), 
            .I1(n4180), .I2(n4597), .I3(\debug_inst/vio0/vio_core_inst/internal_register_select [3]), 
            .O(n4598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77 */ ;
    defparam LUT__10834.LUTMASK = 16'h0f77;
    EFX_LUT4 LUT__10835 (.I0(n4598), .I1(\debug_inst/vio0/vio_core_inst/data_from_biu [1]), 
            .I2(n4182), .O(n4599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c */ ;
    defparam LUT__10835.LUTMASK = 16'h5c5c;
    EFX_LUT4 LUT__10836 (.I0(n4599), .I1(\debug_inst/vio0/vio_core_inst/data_out_shift_reg [2]), 
            .I2(n4185), .O(\debug_inst/vio0/vio_core_inst/n546 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1460)
    defparam LUT__10836.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__10837 (.I0(\debug_inst/vio0/vio_core_inst/word_count [9]), 
            .I1(\debug_inst/vio0/vio_core_inst/word_count [8]), .O(n4600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__10837.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__10838 (.I0(\debug_inst/vio0/vio_core_inst/word_count [12]), 
            .I1(\debug_inst/vio0/vio_core_inst/word_count [11]), .I2(\debug_inst/vio0/vio_core_inst/word_count [10]), 
            .O(n4601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10838.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10839 (.I0(n4158), .I1(n4159), .I2(n4600), .I3(n4601), 
            .O(n4602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10839.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10840 (.I0(\debug_inst/vio0/vio_core_inst/word_count [13]), 
            .I1(n4602), .O(n4603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10840.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10841 (.I0(\debug_inst/vio0/vio_core_inst/word_count [14]), 
            .I1(n4603), .O(n4604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10841.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10842 (.I0(\debug_inst/edb_user_dr [60]), .I1(n4604), 
            .I2(\debug_inst/vio0/vio_core_inst/word_count [15]), .I3(n4139), 
            .O(\debug_inst/vio0/vio_core_inst/data_to_word_counter [15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1438)
    defparam LUT__10842.LUTMASK = 16'haa3c;
    EFX_LUT4 LUT__10843 (.I0(\debug_inst/edb_user_dr [59]), .I1(n4603), 
            .I2(\debug_inst/vio0/vio_core_inst/word_count [14]), .I3(n4139), 
            .O(\debug_inst/vio0/vio_core_inst/data_to_word_counter [14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1438)
    defparam LUT__10843.LUTMASK = 16'haa3c;
    EFX_LUT4 LUT__10844 (.I0(\debug_inst/edb_user_dr [58]), .I1(n4602), 
            .I2(\debug_inst/vio0/vio_core_inst/word_count [13]), .I3(n4139), 
            .O(\debug_inst/vio0/vio_core_inst/data_to_word_counter [13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1438)
    defparam LUT__10844.LUTMASK = 16'haa3c;
    EFX_LUT4 LUT__10845 (.I0(n4160), .I1(n4600), .O(n4605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10845.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10846 (.I0(\debug_inst/vio0/vio_core_inst/word_count [11]), 
            .I1(\debug_inst/vio0/vio_core_inst/word_count [10]), .I2(n4605), 
            .O(n4606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10846.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10847 (.I0(\debug_inst/edb_user_dr [57]), .I1(n4606), 
            .I2(\debug_inst/vio0/vio_core_inst/word_count [12]), .I3(n4139), 
            .O(\debug_inst/vio0/vio_core_inst/data_to_word_counter [12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1438)
    defparam LUT__10847.LUTMASK = 16'haa3c;
    EFX_LUT4 LUT__10848 (.I0(\debug_inst/vio0/vio_core_inst/word_count [10]), 
            .I1(n4605), .I2(\debug_inst/vio0/vio_core_inst/word_count [11]), 
            .O(n4607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b */ ;
    defparam LUT__10848.LUTMASK = 16'h4b4b;
    EFX_LUT4 LUT__10849 (.I0(n4607), .I1(\debug_inst/edb_user_dr [56]), 
            .I2(n4139), .O(\debug_inst/vio0/vio_core_inst/data_to_word_counter [11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1438)
    defparam LUT__10849.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__10850 (.I0(\debug_inst/edb_user_dr [55]), .I1(n4605), 
            .I2(\debug_inst/vio0/vio_core_inst/word_count [10]), .I3(n4139), 
            .O(\debug_inst/vio0/vio_core_inst/data_to_word_counter [10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1438)
    defparam LUT__10850.LUTMASK = 16'haa3c;
    EFX_LUT4 LUT__10851 (.I0(n4605), .I1(n4161), .I2(\debug_inst/edb_user_dr [54]), 
            .I3(n4139), .O(\debug_inst/vio0/vio_core_inst/data_to_word_counter [9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1438)
    defparam LUT__10851.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__10852 (.I0(\debug_inst/edb_user_dr [53]), .I1(n4160), 
            .I2(\debug_inst/vio0/vio_core_inst/word_count [8]), .I3(n4139), 
            .O(\debug_inst/vio0/vio_core_inst/data_to_word_counter [8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1438)
    defparam LUT__10852.LUTMASK = 16'haa3c;
    EFX_LUT4 LUT__10853 (.I0(\debug_inst/vio0/vio_core_inst/word_count [6]), 
            .I1(\debug_inst/vio0/vio_core_inst/word_count [5]), .I2(\debug_inst/vio0/vio_core_inst/word_count [4]), 
            .I3(n4158), .O(n4608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10853.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10854 (.I0(\debug_inst/edb_user_dr [52]), .I1(n4608), 
            .I2(\debug_inst/vio0/vio_core_inst/word_count [7]), .I3(n4139), 
            .O(\debug_inst/vio0/vio_core_inst/data_to_word_counter [7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1438)
    defparam LUT__10854.LUTMASK = 16'haa3c;
    EFX_LUT4 LUT__10855 (.I0(\debug_inst/vio0/vio_core_inst/word_count [5]), 
            .I1(\debug_inst/vio0/vio_core_inst/word_count [4]), .I2(n4158), 
            .I3(\debug_inst/vio0/vio_core_inst/word_count [6]), .O(n4609)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h10ef */ ;
    defparam LUT__10855.LUTMASK = 16'h10ef;
    EFX_LUT4 LUT__10856 (.I0(\debug_inst/edb_user_dr [51]), .I1(n4609), 
            .I2(n4139), .O(\debug_inst/vio0/vio_core_inst/data_to_word_counter [6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1438)
    defparam LUT__10856.LUTMASK = 16'ha3a3;
    EFX_LUT4 LUT__10857 (.I0(\debug_inst/vio0/vio_core_inst/word_count [4]), 
            .I1(n4158), .I2(\debug_inst/vio0/vio_core_inst/word_count [5]), 
            .O(n4610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b */ ;
    defparam LUT__10857.LUTMASK = 16'h4b4b;
    EFX_LUT4 LUT__10858 (.I0(\debug_inst/edb_user_dr [50]), .I1(n4610), 
            .I2(n4139), .O(\debug_inst/vio0/vio_core_inst/data_to_word_counter [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1438)
    defparam LUT__10858.LUTMASK = 16'ha3a3;
    EFX_LUT4 LUT__10859 (.I0(\debug_inst/edb_user_dr [49]), .I1(n4158), 
            .I2(\debug_inst/vio0/vio_core_inst/word_count [4]), .I3(n4139), 
            .O(\debug_inst/vio0/vio_core_inst/data_to_word_counter [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1438)
    defparam LUT__10859.LUTMASK = 16'haa3c;
    EFX_LUT4 LUT__10860 (.I0(\debug_inst/vio0/vio_core_inst/word_count [0]), 
            .I1(\debug_inst/vio0/vio_core_inst/word_count [2]), .I2(\debug_inst/vio0/vio_core_inst/word_count [1]), 
            .I3(\debug_inst/vio0/vio_core_inst/word_count [3]), .O(n4611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h01fe */ ;
    defparam LUT__10860.LUTMASK = 16'h01fe;
    EFX_LUT4 LUT__10861 (.I0(\debug_inst/edb_user_dr [48]), .I1(n4611), 
            .I2(n4139), .O(\debug_inst/vio0/vio_core_inst/data_to_word_counter [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1438)
    defparam LUT__10861.LUTMASK = 16'ha3a3;
    EFX_LUT4 LUT__10862 (.I0(\debug_inst/vio0/vio_core_inst/word_count [0]), 
            .I1(\debug_inst/vio0/vio_core_inst/word_count [1]), .I2(\debug_inst/vio0/vio_core_inst/word_count [2]), 
            .O(n4612)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1e1e */ ;
    defparam LUT__10862.LUTMASK = 16'h1e1e;
    EFX_LUT4 LUT__10863 (.I0(\debug_inst/edb_user_dr [47]), .I1(n4612), 
            .I2(n4139), .O(\debug_inst/vio0/vio_core_inst/data_to_word_counter [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1438)
    defparam LUT__10863.LUTMASK = 16'ha3a3;
    EFX_LUT4 LUT__10864 (.I0(\debug_inst/edb_user_dr [46]), .I1(\debug_inst/vio0/vio_core_inst/word_count [0]), 
            .I2(\debug_inst/vio0/vio_core_inst/word_count [1]), .I3(n4139), 
            .O(\debug_inst/vio0/vio_core_inst/data_to_word_counter [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haac3 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1438)
    defparam LUT__10864.LUTMASK = 16'haac3;
    EFX_LUT4 LUT__10865 (.I0(n4154), .I1(\debug_inst/vio0/vio_core_inst/n408 [5]), 
            .O(\debug_inst/vio0/vio_core_inst/n422 [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1429)
    defparam LUT__10865.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10866 (.I0(n4154), .I1(\debug_inst/vio0/vio_core_inst/n408 [4]), 
            .O(\debug_inst/vio0/vio_core_inst/n422 [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1429)
    defparam LUT__10866.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10867 (.I0(n4154), .I1(\debug_inst/vio0/vio_core_inst/n408 [3]), 
            .O(\debug_inst/vio0/vio_core_inst/n422 [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1429)
    defparam LUT__10867.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10868 (.I0(n4154), .I1(\debug_inst/vio0/vio_core_inst/n408 [2]), 
            .O(\debug_inst/vio0/vio_core_inst/n422 [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1429)
    defparam LUT__10868.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10869 (.I0(n4154), .I1(\debug_inst/vio0/vio_core_inst/n408 [1]), 
            .O(\debug_inst/vio0/vio_core_inst/n422 [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1429)
    defparam LUT__10869.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10896 (.I0(\debug_inst/edb_user_dr [66]), .I1(\debug_inst/vio0/vio_core_inst/incremented_address [5]), 
            .I2(n4139), .O(\debug_inst/vio0/vio_core_inst/data_to_addr_counter [5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1401)
    defparam LUT__10896.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__10897 (.I0(\debug_inst/edb_user_dr [65]), .I1(\debug_inst/vio0/vio_core_inst/incremented_address [4]), 
            .I2(n4139), .O(\debug_inst/vio0/vio_core_inst/data_to_addr_counter [4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1401)
    defparam LUT__10897.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__10898 (.I0(\debug_inst/edb_user_dr [64]), .I1(\debug_inst/vio0/vio_core_inst/incremented_address [3]), 
            .I2(n4139), .O(\debug_inst/vio0/vio_core_inst/data_to_addr_counter [3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1401)
    defparam LUT__10898.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__10899 (.I0(\debug_inst/edb_user_dr [63]), .I1(\debug_inst/vio0/vio_core_inst/incremented_address [2]), 
            .I2(n4139), .O(\debug_inst/vio0/vio_core_inst/data_to_addr_counter [2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1401)
    defparam LUT__10899.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__10900 (.I0(\debug_inst/edb_user_dr [62]), .I1(\debug_inst/vio0/vio_core_inst/incremented_address [1]), 
            .I2(n4139), .O(\debug_inst/vio0/vio_core_inst/data_to_addr_counter [1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1401)
    defparam LUT__10900.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__10901 (.I0(n4217), .I1(\debug_inst/vio0/vio_core_inst/address_counter [1]), 
            .O(n4613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__10901.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__10902 (.I0(n4170), .I1(n4172), .I2(n4173), .I3(n4613), 
            .O(\debug_inst/vio0/vio_core_inst/n2952 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(1866)
    defparam LUT__10902.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10903 (.I0(\debug_inst/vio0/vio_core_inst/module_state [1]), 
            .I1(\debug_inst/vio0/vio_core_inst/module_state [2]), .I2(\debug_inst/vio0/vio_core_inst/module_state [0]), 
            .O(n4614)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__10903.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__10904 (.I0(bscan_SEL), .I1(bscan_UPDATE), .I2(\debug_inst/edb_user_dr [81]), 
            .O(\debug_inst/debug_hub_inst/n265 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(435)
    defparam LUT__10904.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10905 (.I0(n4614), .I1(\debug_inst/vio0/vio_core_inst/module_state [2]), 
            .I2(\debug_inst/vio0/vio_core_inst/module_state [3]), .I3(\debug_inst/debug_hub_inst/n265 ), 
            .O(\debug_inst/debug_hub_inst/n267 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(435)
    defparam LUT__10905.LUTMASK = 16'hc500;
    EFX_LUT4 LUT__10906 (.I0(bscan_SEL), .I1(bscan_SHIFT), .O(\debug_inst/debug_hub_inst/n96 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;   // /home/lalli/Downloads/Efinity_stuff/testing_PLLs/debug_top.v(428)
    defparam LUT__10906.LUTMASK = 16'h8888;
    EFX_GBUFCE CLKBUF__2 (.CE(1'b1), .I(clk_1), .O(\clk_1~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__2.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__1 (.CE(1'b1), .I(clk_0), .O(\clk_0~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__1.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__0 (.CE(1'b1), .I(bscan_TCK), .O(\bscan_TCK~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__0.CE_POLARITY = 1'b1;
    
endmodule

//
// Verific Verilog Description of module EFX_LUT4_f0a24934_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f0a24934_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f0a24934_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f0a24934_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f0a24934_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f0a24934_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f0a24934_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f0a24934_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f0a24934_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_f0a24934_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f0a24934_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE_f0a24934_0
// module not written out since it is a black box. 
//

